CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 130 30 150 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 136 261 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7223 0 0
2
42826.4 0
0
13 Logic Switch~
5 178 261 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3641 0 0
2
42826.4 1
0
13 Logic Switch~
5 258 261 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3104 0 0
2
42826.4 2
0
13 Logic Switch~
5 216 261 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3296 0 0
2
42826.4 3
0
13 Logic Switch~
5 300 261 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8534 0 0
2
42826.4 4
0
13 Logic Switch~
5 294 168 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
949 0 0
2
42826.4 5
0
13 Logic Switch~
5 210 168 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3371 0 0
2
42826.4 6
0
13 Logic Switch~
5 252 168 0 1 11
0 38
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7311 0 0
2
42826.4 7
0
13 Logic Switch~
5 172 168 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
42826.4 8
0
13 Logic Switch~
5 130 168 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3526 0 0
2
42826.4 9
0
8 2-In OR~
219 315 648 0 3 22
0 3 4 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4129 0 0
2
42826.5 1
0
7 74LS283
152 535 462 0 14 29
0 25 24 23 22 2 8 8 2 2
21 20 19 18 13
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
6278 0 0
2
42826.4 3
0
7 Ground~
168 495 522 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3482 0 0
2
42826.4 2
0
7 Ground~
168 675 495 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8323 0 0
2
42826.4 1
0
7 74LS283
152 731 461 0 14 29
0 10 11 12 3 2 2 2 2 13
17 16 15 14 41
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
3984 0 0
2
42826.4 0
0
9 2-In AND~
219 387 495 0 3 22
0 9 7 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7622 0 0
2
42826.4 0
0
12 Hex Display~
7 802 308 0 16 19
10 14 15 16 17 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
816 0 0
2
42826.4 1
0
12 Hex Display~
7 883 308 0 16 19
10 18 19 20 21 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4656 0 0
2
42826.4 0
0
7 Ground~
168 144 675 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6356 0 0
2
42826.4 0
0
6 74LS85
106 225 621 0 14 29
0 25 24 23 22 6 2 2 6 42
43 44 45 46 4
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
3 U10
-10 -62 11 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7479 0 0
2
42826.4 0
0
6 74LS85
106 225 504 0 14 29
0 25 24 23 22 2 2 6 6 47
48 49 27 28 29
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U4
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5690 0 0
2
42826.4 10
0
6 74LS85
106 225 387 0 14 29
0 10 11 12 3 2 2 2 6 27
28 29 9 50 51
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5617 0 0
2
42826.4 9
0
2 +V
167 117 414 0 1 3
0 6
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3903 0 0
2
42826.4 8
0
14 Logic Display~
6 315 387 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4452 0 0
2
42826.4 6
0
7 74LS283
152 490 201 0 14 29
0 40 39 38 37 36 35 34 33 2
25 24 23 22 30
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
6282 0 0
2
42826.4 3
0
7 Ground~
168 450 261 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7187 0 0
2
42826.4 2
0
7 Ground~
168 639 288 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6866 0 0
2
42826.4 1
0
7 74LS283
152 686 200 0 14 29
0 2 2 2 31 2 2 2 32 30
10 11 12 3 52
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
7670 0 0
2
42826.4 0
0
123
5 0 2 0 0 4096 0 22 0 0 74 3
193 396
145 396
145 405
1 -2303 3 0 0 4096 0 11 0 0 3 2
302 639
283 639
-10361022 0 1 0 0 4128 0 0 0 0 0 2
283 615
283 651
14 2 4 0 0 4224 0 20 11 0 0 2
257 657
302 657
0 0 5 0 0 128 0 0 0 0 0 2
351 657
351 657
5 0 6 0 0 4096 0 20 0 0 7 2
193 630
117 630
8 0 6 0 0 8320 0 20 0 0 67 3
193 657
117 657
117 539
0 0 2 0 0 0 0 0 0 9 66 2
180 639
144 639
6 7 2 0 0 0 0 20 20 0 0 4
193 639
180 639
180 648
193 648
0 0 2 0 0 4096 0 0 0 74 66 2
145 414
145 522
2 3 7 0 0 8320 0 16 11 0 0 4
363 504
351 504
351 648
348 648
3 0 8 0 0 4096 0 16 0 0 23 3
408 495
450 495
450 480
1 1 9 0 0 8320 0 16 24 0 0 4
363 486
351 486
351 405
315 405
1 -2300 10 0 0 4224 0 15 0 0 31 2
699 425
661 425
2 -2301 11 0 0 4224 0 15 0 0 31 2
699 434
661 434
3 -2302 12 0 0 4224 0 15 0 0 31 2
699 443
661 443
4 -2303 3 0 0 4224 0 15 0 0 31 2
699 452
661 452
6 0 2 0 0 0 0 15 0 0 21 2
699 470
675 470
7 0 2 0 0 0 0 15 0 0 21 2
699 479
675 479
8 1 2 0 0 0 0 15 14 0 0 3
699 488
699 489
675 489
5 1 2 0 0 0 0 15 14 0 0 3
699 461
675 461
675 489
14 9 13 0 0 8320 0 12 15 0 0 3
567 507
567 506
699 506
7 6 8 0 0 4224 0 12 12 0 0 4
503 480
450 480
450 471
503 471
8 0 2 0 0 0 0 12 0 0 25 2
503 489
496 489
0 5 2 0 0 0 0 0 12 32 0 3
496 507
496 462
503 462
13 -2303 14 0 0 4096 0 15 0 0 30 2
763 479
782 479
12 -2302 15 0 0 4096 0 15 0 0 30 2
763 470
782 470
11 -2301 16 0 0 4096 0 15 0 0 30 2
763 461
782 461
10 -2300 17 0 0 4096 0 15 0 0 30 2
763 452
782 452
-10361020 0 1 0 0 4128 0 0 0 0 0 2
782 436
782 484
-10361022 0 1 0 0 4128 0 0 0 0 0 2
661 405
661 457
9 1 2 0 0 0 0 12 13 0 0 3
503 507
495 507
495 516
13 -2303 18 0 0 4224 0 12 0 0 37 2
567 480
587 480
12 -2302 19 0 0 4224 0 12 0 0 37 2
567 471
587 471
11 -2301 20 0 0 4224 0 12 0 0 37 2
567 462
587 462
10 -2300 21 0 0 4224 0 12 0 0 37 2
567 453
587 453
-10361021 0 1 0 0 32 0 0 0 0 0 2
587 438
587 488
4 -2303 22 0 0 4224 0 12 0 0 42 2
503 453
465 453
3 -2302 23 0 0 4224 0 12 0 0 42 2
503 444
465 444
2 -2301 24 0 0 4224 0 12 0 0 42 2
503 435
465 435
1 -2300 25 0 0 4224 0 12 0 0 42 2
503 426
465 426
-10361023 0 1 0 0 32 0 0 0 0 0 2
465 406
465 458
4 -2300 17 0 0 4224 0 17 0 0 52 2
793 332
793 352
3 -2301 16 0 0 4224 0 17 0 0 52 2
799 332
799 352
2 -2302 15 0 0 4224 0 17 0 0 52 2
805 332
805 352
1 -2303 14 0 0 4224 0 17 0 0 52 2
811 332
811 352
4 -2300 21 0 0 0 0 18 0 0 51 2
874 332
874 352
3 -2301 20 0 0 0 0 18 0 0 51 2
880 332
880 352
2 -2302 19 0 0 0 0 18 0 0 51 2
886 332
886 352
1 -2303 18 0 0 0 0 18 0 0 51 2
892 332
892 352
-10361021 0 1 0 0 32 0 0 0 0 0 2
856 352
903 352
-10361020 0 1 0 0 32 0 0 0 0 0 2
775 352
822 352
0 0 26 0 0 0 0 0 0 0 0 2
180 559
180 559
8 7 6 0 0 0 0 21 21 0 0 4
193 540
180 540
180 531
193 531
1 -2300 25 0 0 0 0 20 0 0 59 2
193 594
172 594
2 -2301 24 0 0 0 0 20 0 0 59 2
193 603
172 603
3 -2302 23 0 0 0 0 20 0 0 59 2
193 612
172 612
4 -2303 22 0 0 0 0 20 0 0 59 2
193 621
172 621
-10361023 0 1 0 0 32 0 0 0 0 0 2
172 574
172 626
0 12 9 0 0 128 0 0 22 61 0 2
299 405
257 405
0 1 9 0 0 0 0 0 24 0 0 2
296 405
315 405
9 12 27 0 0 8320 0 22 21 0 0 4
257 360
289 360
289 522
257 522
10 13 28 0 0 8320 0 22 21 0 0 4
257 369
280 369
280 531
257 531
11 14 29 0 0 8320 0 22 21 0 0 4
257 378
271 378
271 540
257 540
5 0 2 0 0 0 0 21 0 0 66 3
193 513
179 513
179 522
6 1 2 0 0 8320 0 21 19 0 0 3
193 522
144 522
144 669
1 0 6 0 0 128 0 23 0 0 54 3
117 423
117 540
180 540
1 -2300 25 0 0 0 0 21 0 0 72 2
193 477
172 477
2 -2301 24 0 0 0 0 21 0 0 72 2
193 486
172 486
3 -2302 23 0 0 0 0 21 0 0 72 2
193 495
172 495
4 -2303 22 0 0 0 0 21 0 0 72 2
193 504
172 504
-10361023 0 1 0 0 32 0 0 0 0 0 2
172 457
172 509
1 8 6 0 0 0 0 23 22 0 0 2
117 423
193 423
6 7 2 0 0 0 0 22 22 0 0 4
193 405
144 405
144 414
193 414
4 -2303 3 0 0 0 0 22 0 0 79 2
193 387
171 387
3 -2302 12 0 0 0 0 22 0 0 79 2
193 378
171 378
2 -2301 11 0 0 0 0 22 0 0 79 2
193 369
171 369
1 -2300 10 0 0 0 0 22 0 0 79 2
193 360
171 360
-10361022 0 1 0 0 32 0 0 0 0 0 2
171 351
171 392
14 9 30 0 0 8320 0 25 28 0 0 3
522 246
522 245
654 245
5 0 2 0 0 0 0 28 0 0 93 2
654 200
639 200
4 -3452 31 0 0 4096 0 28 0 0 95 2
654 191
616 191
8 -3388 32 0 0 4224 0 28 0 0 94 2
654 227
588 227
0 1 2 0 0 0 0 0 28 93 0 3
639 173
639 164
654 164
13 -2303 3 0 0 0 0 28 0 0 89 2
718 218
737 218
12 -2302 12 0 0 0 0 28 0 0 89 2
718 209
737 209
11 -2301 11 0 0 0 0 28 0 0 89 2
718 200
737 200
10 -2300 10 0 0 0 0 28 0 0 89 2
718 191
737 191
-10361022 0 1 0 0 32 0 0 0 0 0 2
737 175
737 223
7 0 2 0 0 0 0 28 0 0 93 2
654 218
639 218
6 0 2 0 0 0 0 28 0 0 93 2
654 209
639 209
3 0 2 0 0 0 0 28 0 0 93 2
654 182
639 182
2 1 2 0 0 0 0 28 27 0 0 3
654 173
639 173
639 282
-881209461 0 1 0 0 32 0 0 0 0 0 2
588 188
588 234
-881209462 0 1 0 0 32 0 0 0 0 0 2
616 144
616 196
9 1 2 0 0 0 0 25 26 0 0 3
458 246
450 246
450 255
13 -2303 22 0 0 0 0 25 0 0 101 2
522 219
542 219
12 -2302 23 0 0 0 0 25 0 0 101 2
522 210
542 210
11 -2301 24 0 0 0 0 25 0 0 101 2
522 201
542 201
10 -2300 25 0 0 0 0 25 0 0 101 2
522 192
542 192
-10361023 0 1 0 0 32 0 0 0 0 0 2
542 177
542 227
8 -3392 33 0 0 4224 0 25 0 0 106 2
458 228
392 228
7 -3391 34 0 0 4288 0 25 0 0 106 2
458 219
392 219
6 -3390 35 0 0 4224 0 25 0 0 106 2
458 210
392 210
5 -3389 36 0 0 4224 0 25 0 0 106 2
458 201
392 201
-881209461 0 1 0 0 32 0 0 0 0 0 2
392 189
392 235
4 -3456 37 0 0 4096 0 25 0 0 111 2
458 192
420 192
3 -3455 38 0 0 4096 0 25 0 0 111 2
458 183
420 183
2 -3454 39 0 0 4096 0 25 0 0 111 2
458 174
420 174
1 -3453 40 0 0 4096 0 25 0 0 111 2
458 165
420 165
-881209462 0 1 0 0 32 0 0 0 0 0 2
420 145
420 197
1 -3392 33 0 0 0 0 5 0 0 117 2
312 261
312 304
1 -3391 34 0 0 0 0 3 0 0 117 2
270 261
270 304
1 -3390 35 0 0 0 0 4 0 0 117 2
228 261
228 304
1 -3389 36 0 0 0 0 2 0 0 117 2
190 261
190 304
1 -3388 32 0 0 0 0 1 0 0 117 2
148 261
148 304
-881209461 0 1 0 0 4256 0 0 0 0 0 2
115 304
329 304
1 -3456 37 0 0 4224 0 6 0 0 123 2
306 168
306 211
1 -3455 38 0 0 4224 0 8 0 0 123 2
264 168
264 211
1 -3454 39 0 0 4224 0 7 0 0 123 2
222 168
222 211
1 -3453 40 0 0 4224 0 9 0 0 123 2
184 168
184 211
1 -3452 31 0 0 4224 0 10 0 0 123 2
142 168
142 211
-881209462 0 1 0 0 48 0 0 0 0 0 2
109 211
323 211
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
