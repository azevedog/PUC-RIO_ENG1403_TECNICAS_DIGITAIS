CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
56
13 Logic Switch~
5 735 202 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89794e-315 0
0
13 Logic Switch~
5 19 657 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
42821.6 0
0
13 Logic Switch~
5 88 693 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
1 D
-4 -26 3 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
42821.6 1
0
13 Logic Switch~
5 87 656 0 1 11
0 29
0
0 0 21344 180
2 0V
-7 -16 7 -8
1 C
-4 -26 3 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
42821.6 2
0
13 Logic Switch~
5 19 694 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
42821.6 3
0
13 Logic Switch~
5 29 313 0 1 11
0 46
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
42821.6 4
0
13 Logic Switch~
5 33 169 0 1 11
0 47
0
0 0 21344 0
2 0V
-7 -16 7 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
42821.6 5
0
7 Ground~
168 915 273 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
5.89794e-315 0
0
7 Ground~
168 776 490 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.89794e-315 0
0
7 Ground~
168 771 365 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
972 0 0
2
5.89794e-315 0
0
12 Hex Display~
7 1014 249 0 18 19
10 8 7 6 5 0 0 0 0 0
0 0 1 1 1 1 0 1 13
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3472 0 0
2
5.89794e-315 0
0
12 Hex Display~
7 956 251 0 16 19
10 4 3 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9998 0 0
2
5.89794e-315 0
0
7 74LS157
122 820 430 0 14 29
0 20 13 15 2 14 60 61 62 63
2 4 3 64 65
0
0 0 4832 0
7 74LS157
-24 -60 25 -52
3 U10
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89794e-315 0
0
7 74LS157
122 817 307 0 14 29
0 20 9 19 10 18 11 17 12 16
2 8 7 6 5
0
0 0 4832 0
7 74LS157
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.89794e-315 0
0
7 Ground~
168 606 307 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
5.89794e-315 0
0
8 2-In OR~
219 308 1186 0 3 22
0 23 22 21
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
3670 0 0
2
42821.6 6
0
9 3-In AND~
219 216 1214 0 4 22
0 28 27 26 22
0
0 0 608 0
6 74LS11
-21 -28 21 -20
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 10 0
1 U
5616 0 0
2
42821.6 7
0
9 2-In AND~
219 215 1167 0 3 22
0 25 24 23
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9323 0 0
2
42821.6 8
0
14 Logic Display~
6 553 789 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89794e-315 5.26354e-315
0
14 Logic Display~
6 517 789 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89794e-315 5.30499e-315
0
14 Logic Display~
6 480 789 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.89794e-315 5.32571e-315
0
14 Logic Display~
6 439 789 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89794e-315 5.34643e-315
0
8 2-In OR~
219 395 1059 0 3 22
0 39 40 30
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
7876 0 0
2
5.89794e-315 5.3568e-315
0
8 2-In OR~
219 316 1033 0 3 22
0 38 37 39
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U15A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
6369 0 0
2
5.89794e-315 5.36716e-315
0
8 2-In OR~
219 303 922 0 3 22
0 36 35 31
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9172 0 0
2
42821.6 9
0
8 2-In OR~
219 292 764 0 3 22
0 34 33 32
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7100 0 0
2
42821.6 10
0
9 3-In AND~
219 217 1120 0 4 22
0 42 41 24 40
0
0 0 608 0
6 74LS11
-21 -28 21 -20
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 7 0
1 U
3820 0 0
2
42821.6 11
0
9 3-In AND~
219 219 1066 0 4 22
0 28 25 26 37
0
0 0 608 0
6 74LS11
-21 -28 21 -20
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 8 0
1 U
7678 0 0
2
42821.6 12
0
9 2-In AND~
219 218 1013 0 3 22
0 28 29 38
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
961 0 0
2
42821.6 13
0
9 Inverter~
13 86 1003 0 2 22
0 26 24
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U8E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
3178 0 0
2
42821.6 14
0
9 Inverter~
13 87 958 0 2 22
0 29 41
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U8D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
3409 0 0
2
42821.6 15
0
9 3-In AND~
219 206 950 0 4 22
0 42 41 24 35
0
0 0 608 0
6 74LS11
-21 -28 21 -20
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 8 0
1 U
3951 0 0
2
42821.6 16
0
9 Inverter~
13 79 888 0 2 22
0 42 28
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U8C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
8885 0 0
2
42821.6 17
0
9 2-In AND~
219 221 898 0 3 22
0 28 27 36
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3780 0 0
2
42821.6 18
0
9 Inverter~
13 86 836 0 2 22
0 27 25
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U8B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9265 0 0
2
42821.6 19
0
9 3-In AND~
219 208 735 0 4 22
0 42 25 26 34
0
0 0 608 0
6 74LS11
-21 -28 21 -20
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 8 0
1 U
9442 0 0
2
5.89794e-315 5.37752e-315
0
9 2-In AND~
219 211 801 0 3 22
0 42 29 33
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9424 0 0
2
5.89794e-315 5.38788e-315
0
9 2-In XOR~
219 283 526 0 3 22
0 45 44 19
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9968 0 0
2
5.89794e-315 5.39306e-315
0
9 2-In AND~
219 215 479 0 3 22
0 44 45 43
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9281 0 0
2
5.89794e-315 5.39824e-315
0
8 2-In OR~
219 659 332 0 3 22
0 47 46 13
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8464 0 0
2
5.89794e-315 5.41896e-315
0
7 74LS157
122 647 249 0 14 29
0 54 53 52 51 50 49 48 44 45
2 12 11 10 9
0
0 0 4832 0
7 74LS157
-24 -60 25 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
42821.6 20
0
6 74LS83
105 351 427 0 14 29
0 47 53 51 49 46 52 50 48 43
15 16 17 18 14
0
0 0 4832 0
6 74LS83
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3171 0 0
2
5.89794e-315 5.43451e-315
0
14 Logic Display~
6 560 383 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89794e-315 5.4371e-315
0
14 Logic Display~
6 418 385 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
42821.6 21
0
14 Logic Display~
6 529 384 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
42821.6 22
0
14 Logic Display~
6 502 385 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
42821.6 23
0
14 Logic Display~
6 474 385 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
42821.6 24
0
14 Logic Display~
6 447 385 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
42821.6 25
0
14 Logic Display~
6 507 198 0 1 2
10 54
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
42821.6 26
0
14 Logic Display~
6 477 200 0 1 2
10 55
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
42821.6 27
0
14 Logic Display~
6 446 201 0 1 2
10 56
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
42821.6 28
0
6 74LS85
106 332 213 0 14 29
0 47 53 51 49 46 52 50 48 59
58 57 56 55 54
0
0 0 5088 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 1 0 0 0
1 U
4292 0 0
2
5.89794e-315 5.43969e-315
0
7 Ground~
168 269 78 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6118 0 0
2
5.89794e-315 5.44228e-315
0
8 Hex Key~
166 86 250 0 11 12
0 45 48 50 52 0 0 0 0 0
6 54
0
0 0 4640 0
0
4 BCDE
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
34 0 0
2
42821.6 29
0
6 74LS85
106 334 98 0 14 29
0 2 2 2 44 2 2 2 45 66
67 68 59 58 57
0
0 0 5088 0
6 74LS85
-21 -52 21 -44
2 U1
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6357 0 0
2
42821.6 30
0
8 Hex Key~
166 100 121 0 11 12
0 44 49 51 53 0 0 0 0 0
7 55
0
0 0 4640 0
0
4 BCDE
-14 -36 14 -28
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
319 0 0
2
42821.6 31
0
122
2 12 3 0 0 4224 0 12 13 0 0 3
959 275
959 430
852 430
1 11 4 0 0 4224 0 12 13 0 0 3
965 275
965 412
852 412
4 14 5 0 0 8320 0 11 14 0 0 3
1005 273
1005 343
849 343
3 13 6 0 0 8320 0 11 14 0 0 3
1011 273
1011 325
849 325
2 12 7 0 0 8320 0 11 14 0 0 3
1017 273
1017 307
849 307
11 1 8 0 0 4224 0 14 11 0 0 3
849 289
1023 289
1023 273
14 0 9 0 0 8192 0 41 0 0 8 3
679 285
679 288
685 288
0 2 9 0 0 12416 0 0 14 0 0 4
677 288
690 288
690 280
785 280
13 4 10 0 0 12416 0 41 14 0 0 4
679 267
726 267
726 298
785 298
12 6 11 0 0 12416 0 41 14 0 0 4
679 249
707 249
707 316
785 316
11 8 12 0 0 8320 0 41 14 0 0 4
679 231
697 231
697 334
785 334
3 2 13 0 0 8320 0 40 13 0 0 3
692 332
692 403
788 403
4 0 2 0 0 8320 0 13 0 0 23 3
788 421
777 421
777 475
1 4 2 0 0 0 0 8 12 0 0 4
915 267
933 267
933 275
947 275
3 4 2 0 0 0 0 12 12 0 0 2
953 275
947 275
5 0 14 0 0 12416 0 13 0 0 80 5
788 430
760 430
760 479
418 479
418 468
3 0 15 0 0 12416 0 13 0 0 79 5
788 412
753 412
753 467
447 467
447 418
9 0 16 0 0 12416 0 14 0 0 78 5
785 343
717 343
717 457
473 457
473 427
7 0 17 0 0 12416 0 14 0 0 76 4
785 325
727 325
727 436
502 436
5 0 18 0 0 12416 0 14 0 0 77 4
785 307
742 307
742 426
529 426
3 0 19 0 0 12288 0 14 0 0 71 4
785 289
735 289
735 415
560 415
1 0 20 0 0 4096 0 14 0 0 25 2
785 271
753 271
10 1 2 0 0 0 0 13 9 0 0 3
782 475
776 475
776 484
1 10 2 0 0 0 0 10 14 0 0 3
771 359
771 352
779 352
1 1 20 0 0 8320 0 13 1 0 0 4
788 394
753 394
753 202
747 202
10 1 2 0 0 0 0 41 15 0 0 3
609 294
606 294
606 301
1 1 2 0 0 0 0 55 53 0 0 3
302 71
302 72
269 72
1 3 21 0 0 4224 0 19 16 0 0 3
553 807
553 1186
341 1186
2 4 22 0 0 12416 0 16 17 0 0 4
295 1195
281 1195
281 1214
237 1214
1 3 23 0 0 12416 0 16 18 0 0 4
295 1177
277 1177
277 1167
236 1167
0 2 24 0 0 8192 0 0 18 50 0 3
125 1127
125 1176
191 1176
0 1 25 0 0 4096 0 0 18 53 0 3
135 1064
135 1158
191 1158
0 3 26 0 0 4096 0 0 17 36 0 3
171 1075
171 1223
192 1223
0 2 27 0 0 4224 0 0 17 63 0 3
142 907
142 1214
192 1214
0 1 28 0 0 4224 0 0 17 54 0 3
159 1057
159 1205
192 1205
0 3 26 0 0 4224 0 0 28 38 0 3
171 744
171 1075
195 1075
0 0 29 0 0 4096 0 0 0 55 67 2
52 958
52 810
3 0 26 0 0 0 0 36 0 0 60 2
184 744
58 744
1 3 30 0 0 4224 0 20 23 0 0 3
517 807
517 1059
428 1059
1 3 31 0 0 8320 0 21 25 0 0 3
480 807
480 922
336 922
3 1 32 0 0 8320 0 26 22 0 0 5
325 764
379 764
379 827
439 827
439 807
2 3 33 0 0 4224 0 26 37 0 0 4
279 773
241 773
241 801
232 801
1 4 34 0 0 4224 0 26 36 0 0 4
279 755
237 755
237 735
229 735
2 4 35 0 0 12416 0 25 32 0 0 4
290 931
265 931
265 950
227 950
3 1 36 0 0 12416 0 34 25 0 0 4
242 898
263 898
263 913
290 913
4 2 37 0 0 12416 0 28 24 0 0 4
240 1066
260 1066
260 1042
303 1042
1 3 38 0 0 4224 0 24 29 0 0 4
303 1024
257 1024
257 1013
239 1013
3 1 39 0 0 12416 0 24 23 0 0 4
349 1033
362 1033
362 1050
382 1050
2 4 40 0 0 4224 0 23 27 0 0 4
382 1068
305 1068
305 1120
238 1120
0 3 24 0 0 4224 0 0 27 59 0 3
125 1001
125 1129
193 1129
0 2 41 0 0 4224 0 0 27 61 0 3
149 950
149 1120
193 1120
0 1 42 0 0 4224 0 0 27 62 0 3
40 941
40 1111
193 1111
0 2 25 0 0 4224 0 0 28 66 0 3
135 836
135 1066
195 1066
0 1 28 0 0 0 0 0 28 56 0 3
159 1001
159 1057
195 1057
1 2 29 0 0 0 0 31 29 0 0 4
72 958
52 958
52 1022
194 1022
0 1 28 0 0 0 0 0 29 64 0 3
159 889
159 1004
194 1004
1 0 27 0 0 0 0 35 0 0 58 2
71 836
46 836
1 0 27 0 0 0 0 5 0 0 63 3
31 694
46 694
46 873
3 2 24 0 0 0 0 32 30 0 0 4
182 959
125 959
125 1003
107 1003
1 1 26 0 0 0 0 3 30 0 0 4
74 693
58 693
58 1003
71 1003
2 2 41 0 0 0 0 32 31 0 0 3
182 950
108 950
108 958
0 1 42 0 0 0 0 0 32 65 0 3
40 915
40 941
182 941
2 0 27 0 0 0 0 34 0 0 58 3
197 907
46 907
46 869
2 1 28 0 0 0 0 33 34 0 0 4
100 888
120 888
120 889
197 889
0 1 42 0 0 0 0 0 33 69 0 5
40 791
40 915
40 915
40 888
64 888
2 2 25 0 0 0 0 35 36 0 0 4
107 836
140 836
140 735
184 735
1 2 29 0 0 8320 0 4 37 0 0 4
73 656
52 656
52 810
187 810
0 1 42 0 0 0 0 0 37 69 0 3
117 791
117 792
187 792
1 1 42 0 0 0 0 36 2 0 0 6
184 726
117 726
117 791
40 791
40 657
31 657
9 3 43 0 0 12416 0 42 39 0 0 4
319 472
295 472
295 479
236 479
3 1 19 0 0 4224 0 38 43 0 0 3
316 526
560 526
560 401
0 2 44 0 0 8192 0 0 38 75 0 3
132 496
132 535
267 535
0 1 45 0 0 8192 0 0 38 74 0 3
148 514
148 517
267 517
0 2 45 0 0 4096 0 0 39 81 0 5
148 353
148 514
148 514
148 488
191 488
0 1 44 0 0 4096 0 0 39 85 0 5
132 341
132 496
132 496
132 470
191 470
1 12 17 0 0 0 0 46 42 0 0 3
502 403
502 436
383 436
1 13 18 0 0 0 0 45 42 0 0 3
529 402
529 445
383 445
11 1 16 0 0 0 0 42 47 0 0 3
383 427
474 427
474 403
10 1 15 0 0 0 0 42 48 0 0 3
383 418
447 418
447 403
1 14 14 0 0 0 0 44 42 0 0 3
418 403
418 472
383 472
0 0 45 0 0 0 0 0 0 84 105 2
148 353
148 283
0 2 46 0 0 8320 0 0 40 96 0 5
258 427
258 361
629 361
629 341
646 341
0 1 47 0 0 8320 0 0 40 100 0 5
313 391
313 345
618 345
618 323
646 323
9 0 45 0 0 12416 0 41 0 0 0 4
615 285
587 285
587 353
145 353
8 0 44 0 0 12416 0 41 0 0 110 5
615 276
582 276
582 341
131 341
131 145
7 0 48 0 0 12416 0 41 0 0 93 5
615 267
576 267
576 334
271 334
271 454
6 0 49 0 0 12416 0 41 0 0 97 5
615 258
572 258
572 329
277 329
277 418
5 0 50 0 0 12416 0 41 0 0 94 5
615 249
567 249
567 324
283 324
283 445
4 0 51 0 0 12416 0 41 0 0 98 5
615 240
560 240
560 317
288 317
288 409
3 0 52 0 0 12416 0 41 0 0 95 5
615 231
554 231
554 311
294 311
294 436
0 2 53 0 0 8320 0 0 41 99 0 5
300 400
300 307
549 307
549 222
615 222
0 1 54 0 0 12288 0 0 41 111 0 4
507 248
542 248
542 213
615 213
8 0 48 0 0 0 0 42 0 0 104 3
319 454
160 454
160 288
0 7 50 0 0 0 0 0 42 103 0 3
170 293
170 445
319 445
6 0 52 0 0 0 0 42 0 0 102 3
319 436
177 436
177 297
0 5 46 0 0 0 0 0 42 101 0 3
187 313
187 427
319 427
0 4 49 0 0 0 0 0 42 109 0 3
210 153
210 418
319 418
0 3 51 0 0 0 0 0 42 108 0 3
220 156
220 409
319 409
2 0 53 0 0 0 0 42 0 0 107 3
319 400
231 400
231 159
0 1 47 0 0 0 0 0 42 106 0 3
241 169
241 391
319 391
5 1 46 0 0 0 0 52 6 0 0 4
300 222
275 222
275 313
41 313
4 6 52 0 0 0 0 54 52 0 0 5
77 274
77 297
279 297
279 231
300 231
7 3 50 0 0 0 0 52 54 0 0 5
300 240
284 240
284 293
83 293
83 274
2 8 48 0 0 0 0 54 52 0 0 5
89 274
89 288
289 288
289 249
300 249
1 8 45 0 0 0 0 54 55 0 0 5
95 274
95 283
295 283
295 134
302 134
1 1 47 0 0 0 0 52 7 0 0 4
300 186
292 186
292 169
45 169
4 2 53 0 0 0 0 56 52 0 0 5
91 145
91 159
288 159
288 195
300 195
3 3 51 0 0 0 0 52 56 0 0 5
300 204
276 204
276 156
97 156
97 145
4 2 49 0 0 0 0 52 56 0 0 5
300 213
283 213
283 153
103 153
103 145
1 4 44 0 0 0 0 56 55 0 0 4
109 145
276 145
276 98
302 98
1 14 54 0 0 8320 0 49 52 0 0 3
507 216
507 249
364 249
13 1 55 0 0 4224 0 52 50 0 0 3
364 240
477 240
477 218
1 12 56 0 0 8320 0 51 52 0 0 3
446 219
446 231
364 231
14 11 57 0 0 8320 0 55 52 0 0 4
366 134
406 134
406 204
364 204
13 10 58 0 0 8320 0 55 52 0 0 4
366 125
401 125
401 195
364 195
12 9 59 0 0 8320 0 55 52 0 0 4
366 116
396 116
396 186
364 186
3 5 2 0 0 0 0 55 55 0 0 4
302 89
302 108
302 108
302 107
6 5 2 0 0 0 0 55 55 0 0 4
302 116
302 121
302 121
302 107
7 6 2 0 0 0 0 55 55 0 0 4
302 125
302 130
302 130
302 116
1 2 2 0 0 0 0 55 55 0 0 4
302 71
302 86
302 86
302 80
3 2 2 0 0 0 0 55 55 0 0 4
302 89
302 94
302 94
302 80
3 2 2 0 0 0 0 55 55 0 0 4
302 89
302 94
302 94
302 80
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
-7 230 78 254
3 238 67 254
8 NUMERO B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
-3 98 82 122
7 106 71 122
8 NUMERO A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
895 113 1052 137
905 121 1041 137
17 COMPARADOR MOSTRA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
905 132 1038 156
915 140 1027 156
14 O MAIOR NUMERO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
610 119 775 143
620 127 764 143
18 Comparador chave 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
622 141 763 165
632 149 752 165
15 Somador chave 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
11 7 104 31
21 15 93 31
9 QUEST�O 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
11 574 104 598
21 582 93 598
9 QUEST�O 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
