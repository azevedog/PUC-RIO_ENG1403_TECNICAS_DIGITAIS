CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 510 6 120 10
176 80 1278 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 281 649 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 CS1
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3701 0 0
2
42877.7 0
0
13 Logic Switch~
5 331 648 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 WE1
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6316 0 0
2
42877.7 1
0
13 Logic Switch~
5 331 112 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 WE
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8734 0 0
2
5.89801e-315 0
0
13 Logic Switch~
5 281 113 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 CS
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7988 0 0
2
5.89801e-315 5.26354e-315
0
2 +V
167 23 871 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3217 0 0
2
42877.7 0
0
7 Ground~
168 43 894 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3965 0 0
2
42877.7 0
0
12 Hex Display~
7 171 830 0 18 19
10 4 5 6 7 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8239 0 0
2
42877.7 0
0
7 Ground~
168 74 954 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
828 0 0
2
42877.7 0
0
7 Pulser~
4 30 569 0 10 12
0 34 35 36 3 0 0 10 10 4
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6187 0 0
2
42877.7 0
0
7 74LS191
135 105 888 0 14 29
0 2 3 8 2 2 2 2 2 37
38 7 6 5 4
0
0 0 4848 0
7 74LS191
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
7107 0 0
2
42877.7 0
0
12 Hex Display~
7 624 577 0 18 19
10 12 11 10 9 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6433 0 0
2
42877.7 2
0
7 Ground~
168 796 644 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8559 0 0
2
42877.7 3
0
2 +V
167 783 607 0 1 3
0 13
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3674 0 0
2
42877.7 4
0
7 74LS283
152 684 631 0 14 29
0 7 6 5 4 2 2 13 2 2
9 10 11 12 39
0
0 0 4848 180
7 74LS283
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
5697 0 0
2
42877.7 5
0
6 1K RAM
79 304 812 0 20 41
0 40 41 42 43 44 45 7 6 5
4 46 47 48 49 18 17 16 15 19
14
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U4
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
3805 0 0
2
42877.7 6
0
12 Hex Display~
7 393 799 0 18 19
10 15 16 17 18 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
7 RESULT1
-24 -38 25 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5219 0 0
2
42877.7 7
0
7 74LS244
143 497 871 0 18 37
0 50 51 52 53 9 10 11 12 54
55 56 57 18 17 16 15 58 14
0
0 0 4848 180
7 74LS244
-24 -60 25 -52
2 U3
-13 -61 1 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 1 0 0 0
1 U
3795 0 0
2
42877.7 8
0
7 74LS244
143 497 335 0 18 37
0 59 60 61 62 25 26 27 28 63
64 65 66 24 23 22 21 67 20
0
0 0 4848 180
7 74LS244
-24 -60 25 -52
2 U1
-13 -61 1 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 1 0 0 0
1 U
3637 0 0
2
42877.7 9
0
12 Hex Display~
7 393 263 0 16 19
10 21 22 23 24 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
6 RESULT
-21 -38 21 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3226 0 0
2
42877.7 10
0
8 Hex Key~
166 681 110 0 11 12
0 28 27 26 25 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 DATA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6966 0 0
2
5.89801e-315 5.30499e-315
0
8 Hex Key~
166 101 107 0 11 12
0 33 32 31 30 0 0 0 0 0
0 48
0
0 0 4656 0
0
7 ADDRESS
-24 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9796 0 0
2
5.89801e-315 5.32571e-315
0
6 1K RAM
79 304 276 0 20 41
0 68 69 70 71 72 73 30 31 32
33 74 75 76 77 24 23 22 21 29
20
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U2
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
5952 0 0
2
5.89801e-315 5.34643e-315
0
85
4 2 3 0 0 16512 0 9 10 0 0 6
60 569
85 569
85 651
66 651
66 870
73 870
0 -1792 4 0 0 4096 0 0 0 10 56 2
180 924
212 924
0 -1791 5 0 0 4096 0 0 0 9 56 2
173 915
212 915
0 -1790 6 0 0 4096 0 0 0 8 56 2
168 905
212 905
0 -1789 7 0 0 4096 0 0 0 7 56 2
162 897
212 897
1 0 8 0 0 4096 0 5 0 0 11 2
23 880
23 879
11 4 7 0 0 128 0 10 7 0 0 3
137 897
162 897
162 854
3 12 6 0 0 4224 0 7 10 0 0 3
168 854
168 906
137 906
13 2 5 0 0 8320 0 10 7 0 0 3
137 915
174 915
174 854
1 14 4 0 0 4224 0 7 10 0 0 3
180 854
180 924
137 924
3 0 8 0 0 4224 0 10 0 0 0 2
67 879
20 879
1 0 2 0 0 8320 0 10 0 0 14 4
67 861
59 861
59 931
73 931
4 1 2 0 0 128 0 10 6 0 0 4
73 888
42 888
42 888
43 888
8 1 2 0 0 0 0 10 8 0 0 3
73 924
73 948
74 948
7 8 2 0 0 0 0 10 10 0 0 2
73 915
73 924
6 7 2 0 0 0 0 10 10 0 0 2
73 906
73 915
5 6 2 0 0 0 0 10 10 0 0 2
73 897
73 906
0 -1597 9 0 0 4096 0 0 0 22 55 2
615 644
591 644
0 -1598 10 0 0 4096 0 0 0 23 55 2
621 635
591 635
0 -1599 11 0 0 4096 0 0 0 24 55 2
627 626
591 626
0 -1600 12 0 0 4096 0 0 0 25 55 2
633 615
591 615
4 10 9 0 0 4096 0 11 14 0 0 3
615 601
615 644
652 644
3 11 10 0 0 4096 0 11 14 0 0 3
621 601
621 635
652 635
2 12 11 0 0 0 0 11 14 0 0 3
627 601
627 626
652 626
1 13 12 0 0 0 0 11 14 0 0 3
633 601
633 617
652 617
1 -1789 7 0 0 8192 0 14 0 0 30 3
716 671
716 709
770 709
2 -1790 6 0 0 0 0 14 0 0 30 4
716 662
739 662
739 694
770 694
3 -1791 5 0 0 0 0 14 0 0 30 4
716 653
743 653
743 681
770 681
4 -1792 4 0 0 0 0 14 0 0 30 4
716 644
749 644
749 667
770 667
-203315 0 1 0 0 4128 0 0 0 0 0 2
770 646
770 758
0 1 2 0 0 128 0 0 12 33 0 3
733 634
796 634
796 638
9 0 2 0 0 0 0 14 0 0 34 3
716 590
733 590
733 607
5 0 2 0 0 0 0 14 0 0 34 3
716 635
733 635
733 624
8 6 2 0 0 0 0 14 14 0 0 6
716 608
733 608
733 607
733 607
733 626
716 626
7 1 13 0 0 4224 0 14 13 0 0 4
716 617
768 617
768 616
783 616
0 18 14 0 0 8320 0 0 17 50 0 4
354 648
534 648
534 866
529 866
1 0 15 0 0 4096 0 16 0 0 44 2
402 823
402 830
2 0 16 0 0 4096 0 16 0 0 43 2
396 823
396 839
3 0 17 0 0 4096 0 16 0 0 42 2
390 823
390 848
4 0 18 0 0 4096 0 16 0 0 41 2
384 823
384 857
15 13 18 0 0 20608 0 15 17 0 0 6
336 830
345 830
345 824
366 824
366 857
459 857
14 16 17 0 0 4224 0 17 15 0 0 6
459 848
369 848
369 835
342 835
342 839
336 839
15 17 16 0 0 4224 0 17 15 0 0 4
459 839
361 839
361 848
336 848
16 18 15 0 0 4224 0 17 15 0 0 4
459 830
356 830
356 857
336 857
5 -1597 9 0 0 4224 0 17 0 0 55 2
523 857
591 857
6 -1598 10 0 0 4224 0 17 0 0 55 2
523 848
591 848
7 -1599 11 0 0 4224 0 17 0 0 55 2
523 839
591 839
8 -1600 12 0 0 4224 0 17 0 0 55 2
523 830
591 830
1 19 19 0 0 12416 0 1 15 0 0 4
293 649
293 688
342 688
342 776
1 20 14 0 0 0 0 2 15 0 0 4
343 648
355 648
355 785
342 785
7 -1789 7 0 0 4224 0 15 0 0 56 2
272 830
212 830
8 -1790 6 0 0 4224 0 15 0 0 56 2
272 839
212 839
9 -1791 5 0 0 128 0 15 0 0 56 2
272 848
212 848
10 -1792 4 0 0 128 0 15 0 0 56 2
272 857
212 857
-11963432 0 1 0 0 4256 0 0 0 0 0 2
591 983
591 608
-203315 0 1 0 0 32 0 0 0 0 0 2
212 976
212 611
0 18 20 0 0 8320 0 0 18 75 0 4
354 112
534 112
534 330
529 330
1 0 21 0 0 4096 0 19 0 0 65 2
402 287
402 294
2 0 22 0 0 4096 0 19 0 0 64 2
396 287
396 303
3 0 23 0 0 4096 0 19 0 0 63 2
390 287
390 312
4 0 24 0 0 4096 0 19 0 0 62 2
384 287
384 321
15 13 24 0 0 20608 0 22 18 0 0 6
336 294
345 294
345 288
366 288
366 321
459 321
14 16 23 0 0 4224 0 18 22 0 0 6
459 312
369 312
369 299
342 299
342 303
336 303
15 17 22 0 0 4224 0 18 22 0 0 4
459 303
361 303
361 312
336 312
16 18 21 0 0 4224 0 18 22 0 0 4
459 294
356 294
356 321
336 321
5 -1597 25 0 0 4096 0 18 0 0 84 2
523 321
591 321
6 -1598 26 0 0 4096 0 18 0 0 84 2
523 312
591 312
7 -1599 27 0 0 4096 0 18 0 0 84 2
523 303
591 303
8 -1600 28 0 0 4096 0 18 0 0 84 2
523 294
591 294
1 -1600 28 0 0 8320 0 20 0 0 84 3
690 134
690 167
591 167
2 -1599 27 0 0 8320 0 20 0 0 84 3
684 134
684 158
591 158
3 -1598 26 0 0 8320 0 20 0 0 84 3
678 134
678 147
591 147
4 -1597 25 0 0 4224 0 20 0 0 84 2
672 134
591 134
1 19 29 0 0 12416 0 4 22 0 0 4
293 113
293 152
342 152
342 240
1 20 20 0 0 0 0 3 22 0 0 4
343 112
355 112
355 249
342 249
4 -1789 30 0 0 8320 0 21 0 0 85 3
92 131
92 165
212 165
3 -1790 31 0 0 8320 0 21 0 0 85 3
98 131
98 157
212 157
2 -1791 32 0 0 8320 0 21 0 0 85 3
104 131
104 149
212 149
1 -1792 33 0 0 8320 0 21 0 0 85 3
110 131
110 141
212 141
7 -1789 30 0 0 0 0 22 0 0 85 2
272 294
212 294
8 -1790 31 0 0 0 0 22 0 0 85 2
272 303
212 303
9 -1791 32 0 0 0 0 22 0 0 85 2
272 312
212 312
10 -1792 33 0 0 0 0 22 0 0 85 2
272 321
212 321
-13326518 0 1 0 0 32 0 0 0 0 0 2
591 447
591 72
-14101669 0 1 0 0 32 0 0 0 0 0 2
212 440
212 75
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
357 606 448 627
366 613 438 628
9 WRITE = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
359 625 440 646
367 631 431 646
8 READ = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
305 41 386 62
313 47 377 62
8 READ = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
303 20 394 41
312 27 384 42
9 WRITE = 0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
