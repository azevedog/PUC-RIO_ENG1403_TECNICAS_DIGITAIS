CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 300 1 120 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 256
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 378 468 0 1 11
0 18
0
0 0 21104 0
2 0V
-6 -16 8 -8
3 CLK
-9 -17 12 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7419 0 0
2
42891.7 0
0
13 Logic Switch~
5 171 324 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
2 RW
-7 -18 7 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
472 0 0
2
42891.7 0
0
13 Logic Switch~
5 477 513 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
5 CLEAR
-18 9 17 17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4714 0 0
2
42891.6 0
0
8 2-In OR~
219 378 603 0 3 22
0 9 8 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9386 0 0
2
42891.8 0
0
9 2-In AND~
219 324 585 0 3 22
0 7 5 9
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7610 0 0
2
42891.8 1
0
9 2-In AND~
219 324 621 0 3 22
0 6 4 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3482 0 0
2
42891.8 0
0
14 Logic Display~
6 909 702 0 1 2
12 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 EMPTY
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3608 0 0
2
42891.8 0
0
14 Logic Display~
6 909 648 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
4 FULL
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6397 0 0
2
42891.8 0
0
2 +V
167 738 531 0 1 3
0 16
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3967 0 0
2
42891.8 0
0
7 Ground~
168 738 765 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8621 0 0
2
42891.8 0
0
6 74LS85
106 783 585 0 14 29
0 16 16 16 16 15 14 13 12 45
46 47 48 4 10
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U9
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
8901 0 0
2
42891.8 0
0
9 Inverter~
13 243 360 0 2 22
0 7 6
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7385 0 0
2
42891.8 0
0
9 2-In AND~
219 477 369 0 3 22
0 6 18 17
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6519 0 0
2
42891.8 0
0
9 2-In AND~
219 477 477 0 3 22
0 18 7 19
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
552 0 0
2
42891.7 0
0
7 74LS191
135 585 657 0 14 29
0 3 18 20 7 2 2 2 2 49
50 15 14 13 12
0
0 0 4848 0
7 74LS191
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
5551 0 0
2
42891.7 0
0
7 Ground~
168 765 387 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8715 0 0
2
42891.7 0
0
7 74LS157
122 783 450 0 14 29
0 7 21 28 22 27 23 26 24 25
2 32 31 30 29
0
0 0 4848 692
7 74LS157
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
9763 0 0
2
42891.7 0
0
7 Ground~
168 531 720 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8443 0 0
2
42891.7 2
0
7 74LS193
137 585 396 0 14 29
0 17 10 20 2 2 2 2 2 51
52 25 26 27 28
0
0 0 4848 0
2 0V
-7 -51 7 -43
7 ENDADDR
-24 -52 25 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
3719 0 0
2
42891.7 1
0
7 74LS193
137 585 522 0 14 29
0 19 11 20 2 2 2 2 2 53
54 24 23 22 21
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
7 STARTAD
-24 -52 25 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
8671 0 0
2
42891.7 0
0
6 74LS85
106 783 711 0 14 29
0 15 14 13 12 2 2 2 2 55
56 57 58 5 11
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U4
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
7168 0 0
2
42891.7 0
0
7 Ground~
168 855 486 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
49 0 0
2
42891.6 0
0
7 Ground~
168 990 486 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6536 0 0
2
42891.6 0
0
12 Hex Display~
7 1224 459 0 18 19
10 44 43 42 41 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
7 BusDATA
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3931 0 0
2
42891.6 0
0
7 74LS245
64 1053 423 0 18 37
0 2 2 2 2 37 38 39 40 59
60 61 62 41 42 43 44 2 7
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 0 0 0 0
1 U
4390 0 0
2
42891.6 0
0
7 74LS244
143 1053 612 0 18 37
0 33 34 35 36 63 64 65 66 41
42 43 44 67 68 69 70 7 71
0
0 0 4848 0
7 74LS244
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 0 0 0 0
1 U
3242 0 0
2
42891.6 0
0
6 1K RAM
79 918 414 0 20 41
0 2 2 2 2 2 2 29 30 31
32 72 73 74 75 37 38 39 40 2
7
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 0 0 0 0
1 U
6760 0 0
2
42891.6 0
0
8 Hex Key~
166 918 540 0 11 12
0 36 35 34 33 0 0 0 0 0
14 69
0
0 0 4656 0
0
5 INPUT
-17 -34 18 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
5760 0 0
2
42891.6 1
0
127
3 1 3 0 0 4224 0 4 15 0 0 4
411 603
541 603
541 630
547 630
2 -5796881 4 0 0 4224 0 6 0 0 18 2
300 630
164 630
2 -389857796 5 0 0 4224 0 5 0 0 18 2
300 594
164 594
1 0 6 0 0 8320 0 6 0 0 5 3
300 612
269 612
269 360
2 1 6 0 0 0 0 12 13 0 0 2
264 360
453 360
0 1 7 0 0 8192 0 0 12 46 0 4
217 324
216 324
216 360
228 360
1 0 7 0 0 4096 0 5 0 0 45 2
300 576
207 576
2 3 8 0 0 12416 0 4 6 0 0 4
365 612
360 612
360 621
345 621
3 1 9 0 0 4224 0 5 4 0 0 4
345 585
360 585
360 594
365 594
14 -247493649 10 0 0 4096 0 11 0 0 19 2
815 621
863 621
2 -247788297 11 0 0 4224 0 20 0 0 18 2
553 504
164 504
2 -247493649 10 0 0 12416 0 19 0 0 18 4
553 378
495 378
495 405
164 405
14 -247788297 11 0 0 0 0 21 0 0 19 2
815 747
863 747
1 -389857796 5 0 0 0 0 7 0 0 19 2
909 720
863 720
1 -5796881 4 0 0 0 0 8 0 0 19 2
909 666
863 666
13 -389857796 5 0 0 128 0 21 0 0 19 2
815 738
863 738
13 -5796881 4 0 0 128 0 11 0 0 19 2
815 612
863 612
-13531751 0 1 0 0 4128 0 0 0 0 0 2
164 369
164 641
-13531751 0 1 0 0 32 0 0 0 0 0 2
863 594
863 759
8 -155985408 12 0 0 4224 0 11 0 0 47 2
751 621
677 621
7 -155985407 13 0 0 4224 0 11 0 0 47 2
751 612
677 612
6 -155985406 14 0 0 4224 0 11 0 0 47 2
751 603
677 603
5 -155985405 15 0 0 4224 0 11 0 0 47 2
751 594
677 594
1 0 16 0 0 4096 0 11 0 0 28 2
751 558
738 558
2 0 16 0 0 0 0 11 0 0 28 2
751 567
738 567
3 0 16 0 0 0 0 11 0 0 28 2
751 576
738 576
4 0 16 0 0 0 0 11 0 0 28 2
751 585
738 585
1 0 16 0 0 4224 0 9 0 0 0 2
738 540
738 591
8 0 2 0 0 4096 0 21 0 0 33 2
751 747
738 747
7 0 2 0 0 0 0 21 0 0 33 2
751 738
738 738
6 0 2 0 0 0 0 21 0 0 33 2
751 729
738 729
5 0 2 0 0 0 0 21 0 0 33 2
751 720
738 720
1 0 2 0 0 4096 0 10 0 0 0 2
738 759
738 714
1 -155985405 15 0 0 0 0 21 0 0 47 2
751 684
677 684
2 -155985406 14 0 0 0 0 21 0 0 47 2
751 693
677 693
3 -155985407 13 0 0 0 0 21 0 0 47 2
751 702
677 702
3 1 17 0 0 4224 0 13 19 0 0 2
498 369
553 369
2 0 7 0 0 4096 0 14 0 0 45 2
453 486
207 486
0 1 18 0 0 4096 0 0 1 40 0 2
434 468
390 468
1 0 18 0 0 0 0 14 0 0 41 2
453 468
433 468
2 2 18 0 0 8320 0 15 13 0 0 4
553 639
433 639
433 378
453 378
3 1 19 0 0 4224 0 14 20 0 0 4
498 477
549 477
549 495
553 495
4 0 2 0 0 0 0 20 0 0 90 2
553 522
531 522
4 0 2 0 0 0 0 19 0 0 90 2
553 396
531 396
0 4 7 0 0 8336 0 0 15 46 0 3
207 324
207 657
553 657
1 0 7 0 0 4224 0 2 0 0 60 2
183 324
727 324
-14101669 0 1 0 0 4256 0 0 0 0 0 2
677 352
677 736
14 -155985408 12 0 0 128 0 15 0 0 47 2
617 693
677 693
13 -155985407 13 0 0 128 0 15 0 0 47 2
617 684
677 684
12 -155985406 14 0 0 128 0 15 0 0 47 2
617 675
677 675
11 -155985405 15 0 0 128 0 15 0 0 47 2
617 666
677 666
0 1 20 0 0 4096 0 0 3 53 0 4
503 513
488 513
488 513
489 513
3 0 20 0 0 8192 0 19 0 0 54 3
547 387
503 387
503 513
3 3 20 0 0 8320 0 20 15 0 0 4
547 513
503 513
503 648
547 648
8 0 2 0 0 0 0 15 0 0 90 2
553 693
531 693
7 0 2 0 0 0 0 15 0 0 90 2
553 684
531 684
6 0 2 0 0 0 0 15 0 0 90 2
553 675
531 675
5 0 2 0 0 0 0 15 0 0 90 2
553 666
531 666
4 -155985408 12 0 0 128 0 21 0 0 47 2
751 711
677 711
0 1 7 0 0 128 0 0 17 92 0 4
971 324
727 324
727 490
751 490
1 10 2 0 0 0 0 16 17 0 0 4
765 381
765 369
745 369
745 409
2 -640 21 0 0 4224 0 17 0 0 47 2
751 481
677 481
4 -639 22 0 0 4224 0 17 0 0 47 2
751 463
677 463
6 -638 23 0 0 4224 0 17 0 0 47 2
751 445
677 445
8 -637 24 0 0 4224 0 17 0 0 47 2
751 427
677 427
9 -1533 25 0 0 4224 0 17 0 0 47 2
751 418
677 418
7 -1534 26 0 0 4224 0 17 0 0 47 2
751 436
677 436
5 -1535 27 0 0 4224 0 17 0 0 47 2
751 454
677 454
3 -1536 28 0 0 4224 0 17 0 0 47 2
751 472
677 472
14 -640 21 0 0 0 0 20 0 0 47 2
617 558
677 558
13 -639 22 0 0 0 0 20 0 0 47 2
617 549
677 549
12 -638 23 0 0 0 0 20 0 0 47 2
617 540
677 540
11 -637 24 0 0 0 0 20 0 0 47 2
617 531
677 531
11 -1533 25 0 0 0 0 19 0 0 47 2
617 405
677 405
12 -1534 26 0 0 0 0 19 0 0 47 2
617 414
677 414
13 -1535 27 0 0 0 0 19 0 0 47 2
617 423
677 423
14 -1536 28 0 0 0 0 19 0 0 47 2
617 432
677 432
7 14 29 0 0 4224 0 27 17 0 0 4
886 432
837 432
837 418
815 418
8 13 30 0 0 4224 0 27 17 0 0 4
886 441
830 441
830 436
815 436
9 12 31 0 0 4224 0 27 17 0 0 4
886 450
829 450
829 454
815 454
10 11 32 0 0 4224 0 27 17 0 0 4
886 459
837 459
837 472
815 472
8 0 2 0 0 0 0 20 0 0 90 2
553 558
531 558
7 0 2 0 0 0 0 20 0 0 90 2
553 549
531 549
6 0 2 0 0 0 0 20 0 0 90 2
553 540
531 540
5 0 2 0 0 0 0 20 0 0 90 2
553 531
531 531
5 0 2 0 0 0 0 19 0 0 90 2
553 405
531 405
6 0 2 0 0 0 0 19 0 0 90 2
553 414
531 414
7 0 2 0 0 0 0 19 0 0 90 2
553 423
531 423
8 0 2 0 0 0 0 19 0 0 90 2
553 432
531 432
1 0 2 0 0 4224 0 18 0 0 0 2
531 714
531 350
0 17 7 0 0 0 0 0 26 92 0 3
971 385
971 576
1015 576
18 20 7 0 0 0 0 25 27 0 0 6
1085 387
1098 387
1098 324
971 324
971 387
956 387
1 4 33 0 0 4224 0 26 28 0 0 3
1021 585
909 585
909 564
3 2 34 0 0 8320 0 28 26 0 0 3
915 564
915 594
1021 594
2 3 35 0 0 8320 0 28 26 0 0 3
921 564
921 603
1021 603
1 4 36 0 0 8320 0 28 26 0 0 3
927 564
927 612
1021 612
1 0 2 0 0 0 0 27 0 0 103 2
886 378
855 378
2 0 2 0 0 0 0 27 0 0 103 2
886 387
855 387
3 0 2 0 0 0 0 27 0 0 103 2
886 396
855 396
4 0 2 0 0 0 0 27 0 0 103 2
886 405
855 405
5 0 2 0 0 0 0 27 0 0 103 2
886 414
855 414
6 0 2 0 0 0 0 27 0 0 103 2
886 423
855 423
1 0 2 0 0 0 0 22 0 0 0 2
855 480
855 360
4 0 2 0 0 0 0 25 0 0 110 2
1021 423
990 423
3 0 2 0 0 0 0 25 0 0 110 2
1021 414
990 414
2 0 2 0 0 0 0 25 0 0 110 2
1021 405
990 405
1 0 2 0 0 0 0 25 0 0 110 2
1021 396
990 396
17 0 2 0 0 0 0 25 0 0 110 2
1015 387
990 387
19 0 2 0 0 0 0 27 0 0 110 2
956 378
990 378
1 0 2 0 0 0 0 23 0 0 0 2
990 480
990 359
15 5 37 0 0 4224 0 27 25 0 0 2
950 432
1021 432
16 6 38 0 0 4224 0 27 25 0 0 2
950 441
1021 441
17 7 39 0 0 4224 0 27 25 0 0 2
950 450
1021 450
18 8 40 0 0 4224 0 27 25 0 0 2
950 459
1021 459
13 -409765629 41 0 0 4096 0 25 0 0 127 2
1085 432
1133 432
14 -409765630 42 0 0 4096 0 25 0 0 127 2
1085 441
1133 441
15 -409765631 43 0 0 4096 0 25 0 0 127 2
1085 450
1133 450
16 -409765632 44 0 0 4096 0 25 0 0 127 2
1085 459
1133 459
12 -409765632 44 0 0 0 0 26 0 0 127 2
1085 612
1133 612
11 -409765631 43 0 0 0 0 26 0 0 127 2
1085 603
1133 603
10 -409765630 42 0 0 0 0 26 0 0 127 2
1085 594
1133 594
9 -409765629 41 0 0 0 0 26 0 0 127 2
1085 585
1133 585
1 -409765632 44 0 0 8320 0 24 0 0 127 3
1233 483
1233 549
1133 549
2 -409765631 43 0 0 8320 0 24 0 0 127 3
1227 483
1227 531
1133 531
3 -409765630 42 0 0 8320 0 24 0 0 127 3
1221 483
1221 514
1133 514
4 -409765629 41 0 0 8320 0 24 0 0 127 3
1215 483
1215 495
1133 495
-13218332 0 1 0 0 32 0 0 0 0 0 2
1133 349
1133 652
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 147
90 733 643 790
98 739 634 784
147 Esse circuito n�o pode ter um clock muito alto devido ao atraso do 
inversor na entrada "RW". Isso permite a fila pular quando cheia ou 
vazia.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
120 329 207 353
127 334 199 350
9 0 - Write
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
199 655 302 679
206 661 294 677
11 0 - CountUp
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
