CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 140 30 200 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 136 261 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
659 0 0
2
5.89794e-315 0
0
13 Logic Switch~
5 178 261 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3800 0 0
2
5.89794e-315 5.26354e-315
0
13 Logic Switch~
5 258 261 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6792 0 0
2
5.89794e-315 5.30499e-315
0
13 Logic Switch~
5 216 261 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3701 0 0
2
5.89794e-315 5.32571e-315
0
13 Logic Switch~
5 300 261 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6316 0 0
2
5.89794e-315 5.34643e-315
0
13 Logic Switch~
5 294 168 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8734 0 0
2
5.89794e-315 5.3568e-315
0
13 Logic Switch~
5 210 168 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7988 0 0
2
5.89794e-315 5.36716e-315
0
13 Logic Switch~
5 252 168 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3217 0 0
2
5.89794e-315 5.37752e-315
0
13 Logic Switch~
5 172 168 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3965 0 0
2
5.89794e-315 5.38788e-315
0
13 Logic Switch~
5 130 168 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8239 0 0
2
5.89794e-315 5.39306e-315
0
7 Ground~
168 450 567 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
828 0 0
2
42826.5 0
0
7 74LS283
152 488 497 0 14 29
0 7 6 5 4 2 3 3 2 2
11 10 9 8 28
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
6187 0 0
2
42826.5 0
0
12 Hex Display~
7 514 218 0 18 19
10 15 14 13 12 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7107 0 0
2
42826.5 1
0
12 Hex Display~
7 595 218 0 18 19
10 8 9 10 11 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6433 0 0
2
42826.5 0
0
7 74LS283
152 193 381 0 14 29
0 27 26 25 24 23 22 21 20 2
7 6 5 4 29
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
8559 0 0
2
42826.5 6
0
7 Ground~
168 153 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3674 0 0
2
42826.5 5
0
6 74LS85
106 198 513 0 14 29
0 7 6 5 4 19 2 2 19 30
31 32 33 34 3
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
3 U11
-10 -62 11 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5697 0 0
2
42826.5 4
0
2 +V
167 99 504 0 1 3
0 19
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3805 0 0
2
42826.5 3
0
7 Ground~
168 117 567 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5219 0 0
2
42826.5 2
0
7 74LS283
152 389 380 0 14 29
0 2 2 2 17 2 2 2 18 3
12 13 14 15 35
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
3795 0 0
2
42826.5 1
0
7 Ground~
168 342 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3637 0 0
2
42826.5 0
0
80
9 0 2 0 0 4096 0 12 0 0 4 2
456 542
450 542
0 0 3 0 0 4096 0 0 0 5 26 2
413 511
357 511
8 0 2 0 0 0 0 12 0 0 4 2
456 524
450 524
1 5 2 0 0 4096 0 11 12 0 0 3
450 561
450 497
456 497
6 7 3 0 0 0 0 12 12 0 0 4
456 506
413 506
413 515
456 515
4 -2303 4 0 0 4096 0 12 0 0 10 2
456 488
434 488
3 -2302 5 0 0 4096 0 12 0 0 10 2
456 479
434 479
2 -2301 6 0 0 4096 0 12 0 0 10 2
456 470
434 470
1 -2300 7 0 0 4096 0 12 0 0 10 2
456 461
434 461
-10361023 0 1 0 0 4128 0 0 0 0 0 2
434 447
434 495
13 -2303 8 0 0 4096 0 12 0 0 15 2
520 515
539 515
12 -2302 9 0 0 4096 0 12 0 0 15 2
520 506
539 506
11 -2301 10 0 0 4096 0 12 0 0 15 2
520 497
539 497
10 -2300 11 0 0 4096 0 12 0 0 15 2
520 488
539 488
-10361021 0 1 0 0 32 0 0 0 0 0 2
539 472
539 520
4 -2300 12 0 0 4224 0 13 0 0 25 2
505 242
505 262
3 -2301 13 0 0 4224 0 13 0 0 25 2
511 242
511 262
2 -2302 14 0 0 4224 0 13 0 0 25 2
517 242
517 262
1 -2303 15 0 0 4224 0 13 0 0 25 2
523 242
523 262
4 -2300 11 0 0 4224 0 14 0 0 24 2
586 242
586 262
3 -2301 10 0 0 4224 0 14 0 0 24 2
592 242
592 262
2 -2302 9 0 0 4224 0 14 0 0 24 2
598 242
598 262
1 -2303 8 0 0 4224 0 14 0 0 24 2
604 242
604 262
-10361021 0 1 0 0 32 0 0 0 0 0 2
568 262
615 262
-10361022 0 1 0 0 32 0 0 0 0 0 2
487 262
534 262
9 14 3 0 0 8320 0 20 17 0 0 3
357 425
357 549
230 549
0 0 16 0 0 0 0 0 0 0 0 2
342 462
342 462
5 0 2 0 0 0 0 20 0 0 40 2
357 380
342 380
4 -3452 17 0 0 4096 0 20 0 0 42 2
357 371
319 371
8 -3388 18 0 0 4224 0 20 0 0 41 2
357 407
291 407
0 1 2 0 0 0 0 0 20 40 0 3
342 353
342 344
357 344
13 -2303 15 0 0 0 0 20 0 0 36 2
421 398
440 398
12 -2302 14 0 0 0 0 20 0 0 36 2
421 389
440 389
11 -2301 13 0 0 0 0 20 0 0 36 2
421 380
440 380
10 -2300 12 0 0 0 0 20 0 0 36 2
421 371
440 371
-10361022 0 1 0 0 32 0 0 0 0 0 2
440 355
440 403
7 0 2 0 0 0 0 20 0 0 40 2
357 398
342 398
6 0 2 0 0 0 0 20 0 0 40 2
357 389
342 389
3 0 2 0 0 0 0 20 0 0 40 2
357 362
342 362
2 1 2 0 0 8320 0 20 21 0 0 3
357 353
342 353
342 435
-881209461 0 1 0 0 32 0 0 0 0 0 2
291 368
291 414
-881209462 0 1 0 0 4128 0 0 0 0 0 2
319 324
319 376
5 0 19 0 0 4224 0 17 0 0 44 2
166 522
99 522
8 1 19 0 0 0 0 17 18 0 0 3
166 549
99 549
99 513
6 0 2 0 0 0 0 17 0 0 46 3
166 531
117 531
117 540
7 1 2 0 0 0 0 17 19 0 0 3
166 540
117 540
117 561
4 -2303 4 0 0 4224 0 17 0 0 48 2
166 513
137 513
-10361023 0 1 0 0 32 0 0 0 0 0 2
137 474
137 522
3 -2302 5 0 0 4224 0 17 0 0 48 2
166 504
137 504
2 -2301 6 0 0 4224 0 17 0 0 48 2
166 495
137 495
1 -2300 7 0 0 4224 0 17 0 0 48 2
166 486
137 486
1 -636 7 0 0 0 0 17 0 0 48 2
166 486
137 486
9 1 2 0 0 0 0 15 16 0 0 3
161 426
153 426
153 435
13 -2303 4 0 0 0 0 15 0 0 58 2
225 399
245 399
12 -2302 5 0 0 0 0 15 0 0 58 2
225 390
245 390
11 -2301 6 0 0 0 0 15 0 0 58 2
225 381
245 381
10 -2300 7 0 0 0 0 15 0 0 58 2
225 372
245 372
-10361023 0 1 0 0 32 0 0 0 0 0 2
245 357
245 407
8 -3392 20 0 0 4224 0 15 0 0 63 2
161 408
95 408
7 -3391 21 0 0 4288 0 15 0 0 63 2
161 399
95 399
6 -3390 22 0 0 4224 0 15 0 0 63 2
161 390
95 390
5 -3389 23 0 0 4224 0 15 0 0 63 2
161 381
95 381
-881209461 0 1 0 0 32 0 0 0 0 0 2
95 369
95 415
4 -3456 24 0 0 4096 0 15 0 0 68 2
161 372
123 372
3 -3455 25 0 0 4096 0 15 0 0 68 2
161 363
123 363
2 -3454 26 0 0 4096 0 15 0 0 68 2
161 354
123 354
1 -3453 27 0 0 4096 0 15 0 0 68 2
161 345
123 345
-881209462 0 1 0 0 32 0 0 0 0 0 2
123 325
123 377
1 -3392 20 0 0 0 0 5 0 0 74 2
312 261
312 304
1 -3391 21 0 0 0 0 3 0 0 74 2
270 261
270 304
1 -3390 22 0 0 0 0 4 0 0 74 2
228 261
228 304
1 -3389 23 0 0 0 0 2 0 0 74 2
190 261
190 304
1 -3388 18 0 0 0 0 1 0 0 74 2
148 261
148 304
-881209461 0 1 0 0 4256 0 0 0 0 0 2
115 304
329 304
1 -3456 24 0 0 4224 0 6 0 0 80 2
306 168
306 211
1 -3455 25 0 0 4224 0 8 0 0 80 2
264 168
264 211
1 -3454 26 0 0 4224 0 7 0 0 80 2
222 168
222 211
1 -3453 27 0 0 4224 0 9 0 0 80 2
184 168
184 211
1 -3452 17 0 0 4224 0 10 0 0 80 2
142 168
142 211
-881209462 0 1 0 0 32 0 0 0 0 0 2
109 211
323 211
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
