CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 200 5 130 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 864 279 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
2 RW
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9910 0 0
2
5.89805e-315 0
0
13 Logic Switch~
5 252 819 0 1 11
0 50
0
0 0 21104 0
2 0V
-6 -16 8 -8
4 Init
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3834 0 0
2
42906.9 0
0
5 7474~
219 1071 612 0 6 22
0 5 5 7 3 72 6
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U16A
23 -61 51 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
3138 0 0
2
42907 0
0
7 74LS191
135 540 585 0 14 29
0 2 42 3 2 44 45 46 47 73
74 8 9 10 11
0
0 0 4336 0
7 74LS191
-24 -51 25 -43
3 U13
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
5409 0 0
2
42906.9 0
0
7 74LS191
135 540 396 0 14 29
0 2 16 3 2 51 52 49 53 42
75 12 13 14 15
0
0 0 4336 0
7 74LS191
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
983 0 0
2
42906.9 0
0
7 Ground~
168 1035 621 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6652 0 0
2
5.89805e-315 0
0
2 +V
167 1044 531 0 1 3
0 5
0
0 0 53616 0
2 5V
-8 -15 6 -7
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4281 0 0
2
5.89805e-315 0
0
14 Logic Display~
6 1134 558 0 1 2
12 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 MATCH
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6847 0 0
2
5.89805e-315 0
0
6 74LS85
106 990 567 0 14 29
0 17 18 19 20 23 24 25 26 2
5 2 76 7 77
0
0 0 4336 0
6 74LS85
-21 -52 21 -44
3 U14
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6543 0 0
2
5.89805e-315 0
0
7 74LS245
64 990 387 0 18 37
0 78 79 80 81 28 29 30 31 82
83 84 85 17 18 19 20 2 27
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
7168 0 0
2
5.89805e-315 5.34643e-315
0
7 Ground~
168 945 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3828 0 0
2
5.89805e-315 5.32571e-315
0
7 Ground~
168 837 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
955 0 0
2
5.89805e-315 5.30499e-315
0
6 1K RAM
79 882 378 0 20 41
0 2 2 8 9 10 11 12 13 14
15 86 87 88 89 28 29 30 31 2
27
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
7782 0 0
2
5.89805e-315 5.26354e-315
0
8 3-In OR~
219 1161 666 0 4 22
0 6 21 4 16
0
0 0 112 0
4 4075
-14 -24 14 -16
4 U11A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
824 0 0
2
5.89805e-315 0
0
7 Ground~
168 486 783 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6983 0 0
2
5.89805e-315 0
0
14 Logic Display~
6 783 630 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 END
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3185 0 0
2
42906.9 1
0
6 74LS85
106 684 621 0 14 29
0 8 9 10 11 38 39 40 41 90
43 91 92 21 93
0
0 0 4336 0
6 74LS85
-21 -52 21 -44
2 U9
-8 -62 6 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4213 0 0
2
42906.9 3
0
9 Inverter~
13 432 819 0 2 22
0 37 3
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U12B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9765 0 0
2
42906.9 4
0
9 Inverter~
13 396 819 0 2 22
0 50 37
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U12A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8986 0 0
2
42906.9 5
0
7 Pulser~
4 1105 702 0 10 12
0 94 95 4 96 0 0 10 10 1
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3273 0 0
2
42906.9 6
0
6 74LS85
106 684 432 0 14 29
0 12 13 14 15 36 35 34 33 97
98 99 100 43 101
0
0 0 4336 0
6 74LS85
-21 -52 21 -44
3 U10
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5636 0 0
2
42906.9 7
0
12 Quad D Flop~
47 360 765 0 9 19
0 57 56 55 54 26 25 24 23 50
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
2 U7
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
327 0 0
2
42906.9 9
0
8 Hex Key~
166 252 693 0 11 12
0 57 56 55 54 0 0 0 0 0
15 70
0
0 0 4656 0
0
7 toMatch
-20 -34 29 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9233 0 0
2
42906.9 10
0
12 Quad D Flop~
47 360 513 0 9 19
0 64 32 63 62 33 34 35 36 50
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
2 U6
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3875 0 0
2
42906.9 11
0
8 Hex Key~
166 297 450 0 11 12
0 64 32 63 62 0 0 0 0 0
4 52
0
0 0 4656 0
0
6 endAd0
-18 -34 24 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9991 0 0
2
42906.9 12
0
8 Hex Key~
166 252 450 0 11 12
0 61 60 59 58 0 0 0 0 0
1 49
0
0 0 4656 0
0
6 endAd1
-17 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3221 0 0
2
42906.9 13
0
12 Quad D Flop~
47 360 585 0 9 19
0 61 60 59 58 41 40 39 38 50
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
2 U5
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8874 0 0
2
42906.9 14
0
12 Quad D Flop~
47 360 405 0 9 19
0 68 67 66 65 47 46 45 44 50
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
2 U4
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7400 0 0
2
42906.9 15
0
8 Hex Key~
166 252 270 0 11 12
0 68 67 66 65 0 0 0 0 0
0 48
0
0 0 4656 0
0
6 begAd1
-17 -34 25 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3623 0 0
2
42906.9 16
0
8 Hex Key~
166 297 270 0 11 12
0 71 48 70 69 0 0 0 0 0
1 49
0
0 0 4656 0
0
6 BegAd0
-18 -34 24 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3311 0 0
2
42906.9 17
0
12 Quad D Flop~
47 360 333 0 9 19
0 71 48 70 69 53 49 52 51 50
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
2 U3
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5736 0 0
2
42906.9 18
0
12 Hex Display~
7 738 774 0 16 19
10 11 10 9 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 Most
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3143 0 0
2
5.89805e-315 0
0
12 Hex Display~
7 1125 324 0 18 19
10 20 19 18 17 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
6 MemVal
-20 -38 22 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5835 0 0
2
5.89805e-315 5.26354e-315
0
12 Hex Display~
7 792 774 0 18 19
10 15 14 13 12 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 Least
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5108 0 0
2
5.89805e-315 5.30499e-315
0
154
0 4 3 0 0 12416 0 0 3 75 0 5
458 819
460 819
460 872
1071 872
1071 624
3 3 4 0 0 8320 0 20 14 0 0 4
1129 693
1135 693
1135 675
1148 675
0 1 5 0 0 4096 0 0 3 4 0 2
1044 549
1071 549
10 0 5 0 0 0 0 9 0 0 10 2
1022 549
1044 549
0 11 2 0 0 4096 0 0 9 6 0 2
1035 558
1022 558
1 9 2 0 0 4096 0 6 9 0 0 3
1035 615
1035 540
1022 540
1 0 6 0 0 8320 0 14 0 0 8 3
1148 657
1134 657
1134 576
6 1 6 0 0 0 0 3 8 0 0 2
1095 576
1134 576
3 13 7 0 0 4224 0 3 9 0 0 2
1047 594
1022 594
1 2 5 0 0 4224 0 7 3 0 0 3
1044 540
1044 576
1047 576
4 -459375289 8 0 0 4096 0 32 0 0 19 2
729 798
729 844
3 -459375290 9 0 0 4096 0 32 0 0 19 2
735 798
735 844
2 -459375291 10 0 0 4096 0 32 0 0 19 2
741 798
741 844
1 -459375292 11 0 0 4096 0 32 0 0 19 2
747 798
747 844
4 -459375293 12 0 0 4096 0 34 0 0 19 2
783 798
783 844
3 -459375294 13 0 0 4096 0 34 0 0 19 2
789 798
789 844
2 -459375295 14 0 0 4096 0 34 0 0 19 2
795 798
795 844
1 -459375296 15 0 0 4096 0 34 0 0 19 2
801 798
801 844
-13993483 0 1 0 0 4128 0 0 0 0 0 2
622 844
852 844
4 -423679570 16 0 0 4224 0 14 0 0 21 2
1194 666
1253 666
-859887186 0 1 0 0 32 0 0 0 0 0 2
1253 651
1253 699
-423679570 2 16 0 0 128 0 0 5 23 0 4
458 332
504 332
504 378
508 378
-859887186 0 1 0 0 48 0 0 0 0 0 2
458 309
458 357
4 -409765629 17 0 0 4096 0 33 0 0 52 2
1116 348
1071 348
3 -409765630 18 0 0 8192 0 33 0 0 52 3
1122 348
1122 360
1071 360
2 -409765631 19 0 0 8192 0 33 0 0 52 3
1128 348
1128 375
1071 375
1 -409765632 20 0 0 8192 0 33 0 0 52 3
1134 348
1134 387
1071 387
1 2 21 0 0 8320 0 16 14 0 0 3
783 648
783 666
1149 666
0 0 22 0 0 0 0 0 0 0 0 2
737 765
737 765
1 -409765629 17 0 0 4224 0 9 0 0 39 2
958 540
873 540
2 -409765630 18 0 0 4224 0 9 0 0 39 2
958 549
873 549
3 -409765631 19 0 0 4224 0 9 0 0 39 2
958 558
873 558
4 -409765632 20 0 0 4224 0 9 0 0 39 2
958 567
873 567
5 -1684541 23 0 0 4224 0 9 0 0 38 2
958 576
918 576
6 -1684542 24 0 0 4224 0 9 0 0 38 2
958 585
918 585
7 -1684543 25 0 0 4224 0 9 0 0 38 2
958 594
918 594
8 -1684544 26 0 0 4224 0 9 0 0 38 2
958 603
918 603
-694978133 0 1 0 0 32 0 0 0 0 0 2
918 648
918 525
-13218332 0 1 0 0 32 0 0 0 0 0 2
873 516
873 650
20 0 27 0 0 8192 0 13 0 0 41 3
920 351
928 351
928 279
1 18 27 0 0 4224 0 1 10 0 0 4
876 279
1036 279
1036 351
1022 351
17 0 2 0 0 0 0 10 0 0 43 2
952 351
945 351
19 1 2 0 0 8192 0 13 11 0 0 3
920 342
945 342
945 444
15 5 28 0 0 4224 0 13 10 0 0 2
914 396
958 396
16 6 29 0 0 4224 0 13 10 0 0 2
914 405
958 405
17 7 30 0 0 4224 0 13 10 0 0 2
914 414
958 414
18 8 31 0 0 4224 0 13 10 0 0 2
914 423
958 423
13 -409765629 17 0 0 0 0 10 0 0 52 2
1022 396
1071 396
14 -409765630 18 0 0 0 0 10 0 0 52 2
1022 405
1071 405
15 -409765631 19 0 0 0 0 10 0 0 52 2
1022 414
1071 414
16 -409765632 20 0 0 0 0 10 0 0 52 2
1022 423
1071 423
-13218332 0 1 0 0 32 0 0 0 0 0 2
1071 325
1071 432
2 0 2 0 0 0 0 13 0 0 54 2
850 351
837 351
1 1 2 0 0 0 0 12 13 0 0 3
837 444
837 342
850 342
3 -459375289 8 0 0 4096 0 13 0 0 63 2
850 360
793 360
4 -459375290 9 0 0 4096 0 13 0 0 63 2
850 369
793 369
5 -459375291 10 0 0 4096 0 13 0 0 63 2
850 378
793 378
6 -459375292 11 0 0 4096 0 13 0 0 63 2
850 387
793 387
7 -459375293 12 0 0 4096 0 13 0 0 63 2
850 396
793 396
8 -459375294 13 0 0 4096 0 13 0 0 63 2
850 405
793 405
9 -459375295 14 0 0 4096 0 13 0 0 63 2
850 414
793 414
10 -459375296 15 0 0 4096 0 13 0 0 63 2
850 423
793 423
-13993483 0 1 0 0 32 0 0 0 0 0 2
793 306
793 434
8 -1684541 23 0 0 0 0 22 0 0 68 2
384 771
418 771
7 -1684542 24 0 0 0 0 22 0 0 68 2
384 759
418 759
6 -1684543 25 0 0 0 0 22 0 0 68 2
384 747
418 747
5 -1684544 26 0 0 0 0 22 0 0 68 2
384 735
418 735
-694978133 0 1 0 0 32 0 0 0 0 0 2
418 721
418 787
4 0 2 0 0 0 0 5 0 0 73 2
508 396
486 396
4 0 2 0 0 0 0 4 0 0 73 2
508 585
486 585
1 0 2 0 0 0 0 4 0 0 73 2
502 558
486 558
1 0 2 0 0 0 0 5 0 0 73 2
502 369
486 369
1 0 2 0 0 4224 0 15 0 0 0 2
486 777
486 366
3 0 3 0 0 0 0 4 0 0 75 2
502 576
460 576
2 3 3 0 0 128 0 18 5 0 0 4
453 819
460 819
460 387
502 387
2 2 32 0 0 4224 0 24 25 0 0 3
336 495
300 495
300 474
5 -6088256 33 0 0 4096 0 24 0 0 131 2
384 483
419 483
6 -6088255 34 0 0 4096 0 24 0 0 131 2
384 495
419 495
7 -6088254 35 0 0 4096 0 24 0 0 131 2
384 507
419 507
8 -6088253 36 0 0 4096 0 24 0 0 131 2
384 519
419 519
1 2 37 0 0 0 0 18 19 0 0 2
417 819
417 819
8 -6088249 38 0 0 4096 0 27 0 0 131 2
384 591
419 591
7 -6088250 39 0 0 4096 0 27 0 0 131 2
384 579
419 579
6 -6088251 40 0 0 4096 0 27 0 0 131 2
384 567
419 567
5 -6088252 41 0 0 4096 0 27 0 0 131 2
384 555
419 555
9 2 42 0 0 8320 0 5 4 0 0 6
578 387
576 387
576 531
495 531
495 567
508 567
13 1 21 0 0 0 0 17 16 0 0 2
716 648
783 648
13 10 43 0 0 8320 0 21 17 0 0 4
716 459
729 459
729 603
716 603
0 1 8 0 0 0 0 0 17 97 0 2
612 594
652 594
0 2 9 0 0 0 0 0 17 98 0 2
602 603
652 603
0 3 10 0 0 4096 0 0 17 99 0 2
594 612
652 612
0 4 11 0 0 4096 0 0 17 100 0 2
585 621
652 621
8 -6088252 41 0 0 12416 0 17 0 0 131 4
652 657
648 657
648 703
419 703
7 -6088251 40 0 0 12416 0 17 0 0 131 4
652 648
639 648
639 693
419 693
6 -6088250 39 0 0 12416 0 17 0 0 131 4
652 639
631 639
631 684
419 684
5 -6088249 38 0 0 12416 0 17 0 0 131 4
652 630
621 630
621 674
419 674
11 -459375289 8 0 0 12416 0 4 0 0 131 4
572 594
612 594
612 666
419 666
12 -459375290 9 0 0 12416 0 4 0 0 131 4
572 603
603 603
603 657
419 657
13 -459375291 10 0 0 12416 0 4 0 0 131 4
572 612
594 612
594 648
419 648
14 -459375292 11 0 0 12416 0 4 0 0 131 4
572 621
585 621
585 638
419 638
5 -6911353 44 0 0 4288 0 4 0 0 131 2
508 594
419 594
6 -6911354 45 0 0 4224 0 4 0 0 131 2
508 603
419 603
7 -6911355 46 0 0 4224 0 4 0 0 131 2
508 612
419 612
8 -6911356 47 0 0 4224 0 4 0 0 131 2
508 621
419 621
2 2 48 0 0 8320 0 30 31 0 0 3
300 294
300 315
336 315
6 -6911359 49 0 0 4096 0 31 0 0 131 2
384 315
419 315
1 0 50 0 0 4096 0 19 0 0 132 2
381 819
360 819
0 1 12 0 0 0 0 0 21 116 0 2
612 405
652 405
0 2 13 0 0 0 0 0 21 117 0 2
602 414
652 414
0 3 14 0 0 4096 0 0 21 118 0 2
594 423
652 423
0 4 15 0 0 4096 0 0 21 124 0 2
585 432
652 432
8 -6088256 33 0 0 12416 0 21 0 0 131 4
652 468
648 468
648 514
419 514
7 -6088255 34 0 0 12416 0 21 0 0 131 4
652 459
639 459
639 504
419 504
6 -6088254 35 0 0 12416 0 21 0 0 131 4
652 450
631 450
631 495
419 495
5 -6088253 36 0 0 12416 0 21 0 0 131 4
652 441
621 441
621 485
419 485
11 -459375293 12 0 0 12416 0 5 0 0 131 4
572 405
612 405
612 477
419 477
12 -459375294 13 0 0 12416 0 5 0 0 131 4
572 414
603 414
603 468
419 468
13 -459375295 14 0 0 12416 0 5 0 0 131 4
572 423
594 423
594 459
419 459
8 -6911353 44 0 0 0 0 28 0 0 131 2
384 411
419 411
7 -6911354 45 0 0 0 0 28 0 0 131 2
384 399
419 399
6 -6911355 46 0 0 0 0 28 0 0 131 2
384 387
419 387
5 -6911356 47 0 0 0 0 28 0 0 131 2
384 375
419 375
8 -6911357 51 0 0 4096 0 31 0 0 131 2
384 339
419 339
14 -459375296 15 0 0 12416 0 5 0 0 131 4
572 432
585 432
585 449
419 449
5 -6911357 51 0 0 4224 0 5 0 0 131 2
508 405
419 405
6 -6911358 52 0 0 4224 0 5 0 0 131 2
508 414
419 414
7 -6911359 49 0 0 4224 0 5 0 0 131 2
508 423
419 423
8 -6911360 53 0 0 4224 0 5 0 0 131 2
508 432
419 432
7 -6911358 52 0 0 0 0 31 0 0 131 2
384 327
419 327
5 -6911360 53 0 0 0 0 31 0 0 131 2
384 303
419 303
-13993483 0 1 0 0 4256 0 0 0 0 0 2
419 280
419 709
1 9 50 0 0 4096 0 2 22 0 0 3
264 819
360 819
360 801
9 9 50 0 0 4224 0 27 22 0 0 2
360 621
360 801
4 4 54 0 0 8320 0 23 22 0 0 3
243 717
243 771
336 771
3 3 55 0 0 4224 0 22 23 0 0 3
336 759
249 759
249 717
2 2 56 0 0 8320 0 23 22 0 0 3
255 717
255 747
336 747
1 1 57 0 0 8320 0 23 22 0 0 3
261 717
261 735
336 735
9 9 50 0 0 0 0 28 24 0 0 2
360 441
360 549
4 4 58 0 0 4224 0 26 27 0 0 3
243 474
243 591
336 591
3 3 59 0 0 8320 0 27 26 0 0 3
336 579
249 579
249 474
2 2 60 0 0 4224 0 26 27 0 0 3
255 474
255 567
336 567
1 1 61 0 0 4224 0 26 27 0 0 3
261 474
261 555
336 555
9 9 50 0 0 0 0 24 27 0 0 2
360 549
360 621
4 4 62 0 0 4224 0 24 25 0 0 3
336 519
288 519
288 474
3 3 63 0 0 4224 0 24 25 0 0 3
336 507
294 507
294 474
1 1 64 0 0 4224 0 24 25 0 0 3
336 483
306 483
306 474
4 4 65 0 0 4224 0 29 28 0 0 3
243 294
243 411
336 411
3 3 66 0 0 8320 0 28 29 0 0 3
336 399
249 399
249 294
2 2 67 0 0 4224 0 29 28 0 0 3
255 294
255 387
336 387
1 1 68 0 0 4224 0 29 28 0 0 3
261 294
261 375
336 375
9 9 50 0 0 0 0 31 28 0 0 2
360 369
360 441
4 4 69 0 0 4224 0 31 30 0 0 3
336 339
288 339
288 294
3 3 70 0 0 4224 0 31 30 0 0 3
336 327
294 327
294 294
1 1 71 0 0 4224 0 31 30 0 0 3
336 303
306 303
306 294
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
250 202 365 223
259 209 355 224
12 Input Params
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
823 224 912 248
831 231 903 247
9 Write = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
670 703 863 727
678 709 854 725
22 Current Memory Address
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
