CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
280 20 1 170 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 558 207 0 1 11
0 10
0
0 0 21088 0
2 0V
-6 -16 8 -8
5 Clear
-22 -15 13 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89803e-315 0
0
13 Logic Switch~
5 306 270 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21216 0
2 5V
-28 -4 -14 4
7 PushPul
-23 9 26 17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89803e-315 0
0
13 Logic Switch~
5 477 261 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21216 0
2 5V
-6 -16 8 -8
3 CLK
-14 -15 7 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89803e-315 0
0
14 Logic Display~
6 450 135 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
4 Full
8 -11 36 -3
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.89803e-315 0
0
14 Logic Display~
6 432 135 0 1 2
12 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 Empty
-42 -10 -7 -2
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89803e-315 0
0
7 Ground~
168 837 333 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
5.89803e-315 0
0
8 Hex Key~
166 846 405 0 11 12
0 23 22 21 20 0 0 0 0 0
15 70
0
0 0 4640 0
0
5 Input
-17 -34 18 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8901 0 0
2
5.89803e-315 5.26354e-315
0
9 2-In AND~
219 405 198 0 3 22
0 9 11 8
0
0 0 96 692
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7361 0 0
2
5.89803e-315 0
0
9 2-In NOR~
219 468 216 0 3 22
0 8 7 12
0
0 0 96 0
6 74LS02
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4747 0 0
2
5.89803e-315 0
0
9 2-In AND~
219 405 234 0 3 22
0 13 11 7
0
0 0 96 692
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
972 0 0
2
5.89803e-315 0
0
9 Inverter~
13 360 243 0 2 22
0 9 13
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3472 0 0
2
5.89803e-315 0
0
9 2-In AND~
219 531 252 0 3 22
0 15 12 14
0
0 0 96 692
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9998 0 0
2
5.89803e-315 0
0
7 74LS191
135 648 270 0 14 29
0 2 14 10 9 2 2 2 2 28
11 16 17 18 19
0
0 0 4832 0
7 74LS191
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89803e-315 5.30499e-315
0
7 Ground~
168 576 324 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89803e-315 0
0
6 1K RAM
79 783 261 0 20 41
0 2 2 2 2 2 2 16 17 18
19 2 2 2 2 24 25 26 27 2
9
0
0 0 4832 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.89803e-315 5.38788e-315
0
7 Ground~
168 738 333 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
5.89803e-315 5.36716e-315
0
7 74LS245
64 900 270 0 18 37
0 29 30 31 32 24 25 26 27 33
34 35 36 6 5 4 3 2 9
0
0 0 4832 0
7 74LS245
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
5.89803e-315 5.3568e-315
0
12 Hex Display~
7 1026 333 0 18 19
10 3 4 5 6 0 0 0 0 0
0 0 1 1 1 1 0 1 13
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
7 BusData
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9323 0 0
2
5.89803e-315 5.32571e-315
0
7 74LS244
143 900 477 0 18 37
0 20 21 22 23 37 38 39 40 6
5 4 3 41 42 43 44 9 45
0
0 0 4832 0
7 74LS244
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
5.89803e-315 5.30499e-315
0
60
12 -409765632 3 0 0 4096 0 19 0 0 13 2
932 477
972 477
11 -409765631 4 0 0 4096 0 19 0 0 13 2
932 468
972 468
10 -409765630 5 0 0 4096 0 19 0 0 13 2
932 459
972 459
9 -409765629 6 0 0 4096 0 19 0 0 13 2
932 450
972 450
1 -409765632 3 0 0 4224 0 18 0 0 13 3
1035 357
1035 423
972 423
2 -409765631 4 0 0 8320 0 18 0 0 13 3
1029 357
1029 405
972 405
3 -409765630 5 0 0 8320 0 18 0 0 13 3
1023 357
1023 386
972 386
4 -409765629 6 0 0 8320 0 18 0 0 13 3
1017 357
1017 369
972 369
13 -409765629 6 0 0 0 0 17 0 0 13 2
932 279
972 279
14 -409765630 5 0 0 0 0 17 0 0 13 2
932 288
972 288
15 -409765631 4 0 0 0 0 17 0 0 13 2
932 297
972 297
16 -409765632 3 0 0 0 0 17 0 0 13 2
932 306
972 306
-13218332 0 1 0 0 4256 0 0 0 0 0 2
972 214
972 486
1 2 7 0 0 4224 0 4 9 0 0 3
450 153
450 225
455 225
1 0 8 0 0 4224 0 5 0 0 30 2
432 153
432 198
17 0 2 0 0 4096 0 17 0 0 22 2
862 234
837 234
17 0 9 0 0 4096 0 19 0 0 24 2
862 441
772 441
14 0 2 0 0 0 0 15 0 0 22 2
815 270
837 270
13 0 2 0 0 0 0 15 0 0 22 2
815 261
837 261
12 0 2 0 0 0 0 15 0 0 22 2
815 252
837 252
11 0 2 0 0 0 0 15 0 0 22 2
815 243
837 243
19 1 2 0 0 8320 0 15 6 0 0 3
821 225
837 225
837 327
20 0 9 0 0 8192 0 15 0 0 25 3
821 234
829 234
829 116
0 0 9 0 0 4096 0 0 0 25 0 3
712 116
712 441
777 441
0 18 9 0 0 8320 0 0 17 32 0 5
334 207
334 116
946 116
946 234
932 234
3 1 10 0 0 8320 0 13 1 0 0 4
610 261
593 261
593 207
570 207
2 0 11 0 0 4096 0 8 0 0 28 2
381 189
370 189
10 2 11 0 0 12416 0 13 10 0 0 6
680 270
694 270
694 172
370 172
370 225
381 225
3 2 7 0 0 0 0 10 9 0 0 4
426 234
432 234
432 225
455 225
1 3 8 0 0 0 0 9 8 0 0 4
455 207
432 207
432 198
426 198
3 2 12 0 0 4224 0 9 12 0 0 2
507 216
507 243
1 1 9 0 0 0 0 8 11 0 0 4
381 207
334 207
334 243
345 243
1 2 13 0 0 4224 0 10 11 0 0 4
381 243
377 243
377 243
381 243
1 0 9 0 0 0 0 11 0 0 41 3
345 243
334 243
334 270
2 3 14 0 0 4224 0 13 12 0 0 2
616 252
552 252
1 1 15 0 0 4224 0 3 12 0 0 2
489 261
507 261
8 0 2 0 0 0 0 13 0 0 46 2
616 306
576 306
7 0 2 0 0 0 0 13 0 0 46 2
616 297
576 297
6 0 2 0 0 0 0 13 0 0 46 2
616 288
576 288
5 0 2 0 0 0 0 13 0 0 46 2
616 279
576 279
1 4 9 0 0 0 0 2 13 0 0 2
318 270
616 270
11 7 16 0 0 4224 0 13 15 0 0 2
680 279
751 279
12 8 17 0 0 4224 0 13 15 0 0 2
680 288
751 288
13 9 18 0 0 4224 0 13 15 0 0 2
680 297
751 297
14 10 19 0 0 4224 0 13 15 0 0 2
680 306
751 306
1 1 2 0 0 0 0 14 13 0 0 3
576 318
576 243
610 243
4 1 20 0 0 8320 0 7 19 0 0 3
837 429
837 450
868 450
3 2 21 0 0 4224 0 7 19 0 0 3
843 429
843 459
868 459
2 3 22 0 0 4224 0 7 19 0 0 3
849 429
849 468
868 468
1 4 23 0 0 4224 0 7 19 0 0 3
855 429
855 477
868 477
15 5 24 0 0 4224 0 15 17 0 0 2
815 279
868 279
16 6 25 0 0 4224 0 15 17 0 0 2
815 288
868 288
17 7 26 0 0 4224 0 15 17 0 0 2
815 297
868 297
18 8 27 0 0 4224 0 15 17 0 0 2
815 306
868 306
6 0 2 0 0 0 0 15 0 0 60 2
751 270
737 270
5 0 2 0 0 0 0 15 0 0 60 2
751 261
737 261
4 0 2 0 0 0 0 15 0 0 60 2
751 252
737 252
3 0 2 0 0 0 0 15 0 0 60 2
751 243
737 243
2 0 2 0 0 0 0 15 0 0 60 2
751 234
737 234
1 1 2 0 0 0 0 15 16 0 0 4
751 225
737 225
737 327
738 327
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 150
453 28 834 112
459 33 827 97
150 Esse circuito n�o pode ter um clock muito alto 
devido ao atraso do inversor na entrada "RW". 
Isso permite a fila pular quando cheia ou 
vazia.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
357 270 546 294
363 275 539 291
22 Push = 0V -> Pull = 5V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
349 286 546 310
355 291 539 307
23 Write = 0V -> Read = 5V
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
