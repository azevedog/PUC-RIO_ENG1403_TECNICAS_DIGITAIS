CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 140 30 50 10
1017 88 1677 988
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1185 184 1298 281
110100498 256
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 18 288 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 X1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8324 0 0
2
42877.6 2
0
13 Logic Switch~
5 17 328 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 X0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3445 0 0
2
42877.6 1
0
13 Logic Switch~
5 611 184 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 CLK
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7543 0 0
2
42877.6 0
0
5 7415~
219 880 468 0 4 22
0 5 4 6 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 4 0
1 U
6187 0 0
2
42877.6 5
0
5 7415~
219 882 522 0 4 22
0 7 4 6 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
5476 0 0
2
42877.6 4
0
14 Logic Display~
6 963 216 0 1 2
12 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Abriu
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3936 0 0
2
42877.6 3
0
14 Logic Display~
6 918 216 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 Travou
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5770 0 0
2
42877.6 2
0
7 Ground~
168 999 594 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7884 0 0
2
42877.6 1
0
12 Hex Display~
7 1026 558 0 18 19
10 3 4 5 2 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3690 0 0
2
42877.6 0
0
6 JK RN~
219 678 324 0 6 22
0 17 15 19 19 6 3
0
0 0 4720 0
7 74LS107
-25 -42 24 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 1 12 4 13 2 3 1 12 4
13 2 3 8 9 11 10 6 5 0
65 0 0 0 2 1 2 0
1 U
3611 0 0
2
42877.6 3
0
2 +V
167 637 351 0 1 3
0 19
0
0 0 61680 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7912 0 0
2
42877.6 2
0
8 2-In OR~
219 603 306 0 3 22
0 16 7 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6416 0 0
2
42877.6 1
0
5 7415~
219 549 297 0 4 22
0 14 11 10 16
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 4 0
1 U
7278 0 0
2
42877.6 0
0
6 JK RN~
219 679 747 0 6 22
0 20 15 21 26 7 5
0
0 0 4720 0
7 74LS107
-25 -42 24 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 1 12 4 13 2 3 1 12 4
13 2 3 8 9 11 10 6 5 0
65 0 0 0 2 1 3 0
1 U
6804 0 0
2
42877.6 7
0
2 +V
167 630 774 0 1 3
0 26
0
0 0 61680 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9568 0 0
2
42877.6 6
0
9 2-In AND~
219 504 711 0 3 22
0 3 13 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
7178 0 0
2
42877.6 5
0
8 2-In OR~
219 540 720 0 3 22
0 24 23 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7982 0 0
2
42877.6 4
0
8 2-In OR~
219 585 729 0 3 22
0 25 22 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
513 0 0
2
42877.6 3
0
9 2-In AND~
219 549 773 0 3 22
0 3 10 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
8190 0 0
2
42877.6 2
0
9 2-In AND~
219 504 744 0 3 22
0 4 3 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
5209 0 0
2
42877.6 1
0
5 7415~
219 603 810 0 4 22
0 3 11 34 21
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 512 3 2 5 0
1 U
7239 0 0
2
42877.6 0
0
6 JK RN~
219 676 549 0 6 22
0 28 15 27 33 14 4
0
0 0 4720 0
7 74LS107
-25 -42 24 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 6 5 1 12 4
13 2 3 8 9 11 10 6 5 0
65 0 0 0 2 2 2 0
1 U
9474 0 0
2
42877.6 8
0
2 +V
167 648 567 0 1 3
0 33
0
0 0 61680 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3783 0 0
2
42877.6 7
0
8 2-In OR~
219 612 531 0 3 22
0 32 29 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
5422 0 0
2
42877.6 6
0
8 2-In OR~
219 567 522 0 3 22
0 31 30 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
8527 0 0
2
42877.6 5
0
9 2-In AND~
219 531 513 0 3 22
0 6 13 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
761 0 0
2
42877.6 4
0
9 2-In AND~
219 531 546 0 3 22
0 11 12 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
7323 0 0
2
42877.6 3
0
9 2-In AND~
219 576 575 0 3 22
0 5 3 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
8543 0 0
2
42877.6 2
0
8 2-In OR~
219 621 621 0 3 22
0 35 3 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 6 0
1 U
4240 0 0
2
42877.6 1
0
5 7415~
219 594 612 0 4 22
0 7 11 10 36
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 512 3 1 5 0
1 U
7857 0 0
2
42877.6 0
0
9 Inverter~
13 153 355 0 2 22
0 10 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
7255 0 0
2
42877.6 0
0
9 Inverter~
13 153 303 0 2 22
0 11 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
7736 0 0
2
42877.6 0
0
7 Ground~
168 63 216 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5435 0 0
2
42877.6 3
0
12 Hex Display~
7 90 180 0 18 19
10 10 11 2 2 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3446 0 0
2
42877.6 0
0
83
1 -256 3 0 0 4112 0 9 0 0 4 2
1035 582
1035 637
2 -255 4 0 0 4112 0 9 0 0 4 2
1029 582
1029 637
3 -254 5 0 0 4112 0 9 0 0 4 2
1023 582
1023 637
-160201 0 1 0 0 4144 0 0 0 0 0 2
943 637
1081 637
3 -57600 6 0 0 4112 0 5 0 0 11 2
858 531
814 531
2 -255 4 0 0 16 0 5 0 0 11 2
858 522
814 522
1 -57598 7 0 0 4112 0 5 0 0 11 2
858 513
814 513
3 -57600 6 0 0 16 0 4 0 0 11 2
856 477
814 477
2 -255 4 0 0 16 0 4 0 0 11 2
856 468
814 468
1 -254 5 0 0 16 0 4 0 0 11 2
856 459
814 459
-160201 0 1 0 0 48 0 0 0 0 0 2
814 436
814 552
4 1 2 0 0 8336 0 9 8 0 0 3
1017 582
1017 588
999 588
1 4 8 0 0 4240 0 7 4 0 0 3
918 234
918 468
901 468
4 1 9 0 0 8336 0 5 6 0 0 3
903 522
963 522
963 234
2 -320 10 0 0 4096 0 19 0 0 47 2
525 782
417 782
5 -57600 6 0 0 0 0 10 0 0 57 2
708 325
735 325
1 0 11 0 0 4096 0 32 0 0 20 3
138 303
93 303
93 288
1 0 10 0 0 0 0 31 0 0 19 3
138 355
99 355
99 328
0 -320 10 0 0 0 0 0 0 83 45 2
99 328
197 328
0 -319 11 0 0 4096 0 0 0 82 45 2
92 288
197 288
0 -57664 12 0 0 4224 0 0 0 0 47 2
585 819
417 819
2 -319 11 0 0 4224 0 21 0 0 47 2
579 810
417 810
1 -256 3 0 0 4096 0 21 0 0 46 2
579 801
335 801
1 -256 3 0 0 0 0 19 0 0 46 2
525 764
335 764
2 -256 3 0 0 0 0 20 0 0 46 2
480 753
335 753
1 -255 4 0 0 4224 0 20 0 0 46 2
480 735
335 735
2 -57663 13 0 0 4096 0 16 0 0 47 2
480 720
417 720
1 -256 3 0 0 0 0 16 0 0 46 4
480 702
338 702
338 708
335 708
3 -320 10 0 0 4224 0 30 0 0 49 4
570 621
411 621
411 620
408 620
2 -319 11 0 0 0 0 30 0 0 49 2
570 612
408 612
1 -57598 7 0 0 4224 0 30 0 0 48 2
570 603
326 603
2 -256 3 0 0 4224 0 29 0 0 48 4
608 630
343 630
343 620
326 620
2 -256 3 0 0 0 0 28 0 0 48 2
552 584
326 584
1 -254 5 0 0 4224 0 28 0 0 48 2
552 566
326 566
2 -57664 12 0 0 0 0 27 0 0 49 2
507 555
408 555
1 -319 11 0 0 0 0 27 0 0 49 2
507 537
408 537
2 -57663 13 0 0 4224 0 26 0 0 49 2
507 522
408 522
1 -57600 6 0 0 4224 0 26 0 0 48 2
507 504
326 504
3 -320 10 0 0 0 0 13 0 0 51 2
525 306
462 306
2 -319 11 0 0 0 0 13 0 0 51 2
525 297
462 297
1 -57599 14 0 0 4224 0 13 0 0 50 2
525 288
380 288
2 -57598 7 0 0 0 0 12 0 0 50 2
590 315
380 315
2 -57664 12 0 0 0 0 31 0 0 45 2
174 355
197 355
2 -57663 13 0 0 0 0 32 0 0 45 2
174 303
197 303
-2895 0 1 0 0 32 0 0 0 0 0 2
197 260
197 390
-160201 0 1 0 0 32 0 0 0 0 0 2
335 697
335 831
-2895 0 1 0 0 32 0 0 0 0 0 2
417 693
417 830
-160201 0 1 0 0 32 0 0 0 0 0 2
326 490
326 624
-2895 0 1 0 0 32 0 0 0 0 0 2
408 486
408 623
-160201 0 1 0 0 32 0 0 0 0 0 2
380 247
380 381
-2895 0 1 0 0 32 0 0 0 0 0 2
462 243
462 380
5 -57598 7 0 0 128 0 14 0 0 57 2
709 748
735 748
6 -254 5 0 0 128 0 14 0 0 57 2
703 730
735 730
5 -57599 14 0 0 128 0 22 0 0 57 2
706 550
735 550
6 -255 4 0 0 128 0 22 0 0 57 2
700 532
735 532
6 -256 3 0 0 128 0 10 0 0 57 2
702 307
735 307
-160201 0 1 0 0 4256 0 0 0 0 0 2
735 256
735 827
2 2 15 0 0 8192 0 22 14 0 0 3
645 541
648 541
648 739
2 2 15 0 0 8320 0 10 22 0 0 3
647 316
645 316
645 541
1 2 15 0 0 0 0 3 10 0 0 3
623 184
647 184
647 316
4 1 16 0 0 4224 0 13 12 0 0 2
570 297
590 297
3 1 17 0 0 8320 0 12 10 0 0 3
636 306
636 307
654 307
0 0 18 0 0 0 0 0 0 0 0 2
700 363
700 363
4 0 19 0 0 8192 0 10 0 0 65 3
678 355
678 363
654 363
1 3 19 0 0 12416 0 11 10 0 0 4
637 360
637 363
654 363
654 325
3 1 20 0 0 8320 0 18 14 0 0 3
618 729
618 730
655 730
3 4 21 0 0 4224 0 14 21 0 0 3
655 748
655 810
624 810
2 3 22 0 0 8320 0 18 19 0 0 3
572 738
570 738
570 773
2 3 23 0 0 8320 0 17 20 0 0 3
527 729
525 729
525 744
1 3 24 0 0 4224 0 17 16 0 0 2
527 711
525 711
1 3 25 0 0 4224 0 18 17 0 0 2
572 720
573 720
1 4 26 0 0 12416 0 15 14 0 0 5
630 783
631 783
631 785
679 785
679 778
3 3 27 0 0 16512 0 29 22 0 0 6
654 621
664 621
664 593
631 593
631 550
652 550
3 1 28 0 0 8320 0 24 22 0 0 3
645 531
645 532
652 532
2 3 29 0 0 8320 0 24 28 0 0 3
599 540
597 540
597 575
2 3 30 0 0 8320 0 25 27 0 0 3
554 531
552 531
552 546
3 1 31 0 0 4224 0 26 25 0 0 2
552 513
554 513
3 1 32 0 0 4224 0 25 24 0 0 2
600 522
599 522
1 4 33 0 0 8320 0 23 22 0 0 4
648 576
648 586
676 586
676 580
3 0 2 0 0 0 0 34 0 0 81 3
87 204
87 210
81 210
4 1 2 0 0 128 0 34 33 0 0 3
81 204
81 210
63 210
1 2 11 0 0 128 0 1 34 0 0 3
30 288
93 288
93 204
1 1 10 0 0 128 0 2 34 0 0 3
29 328
99 328
99 204
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
