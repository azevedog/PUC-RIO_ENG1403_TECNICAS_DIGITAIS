CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 0 8 150 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.585492 0.500000
176 80 1278 659
42991634 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 517 633 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9953 0 0
2
5.89796e-315 5.34643e-315
0
13 Logic Switch~
5 510 679 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
361 0 0
2
5.89796e-315 5.32571e-315
0
13 Logic Switch~
5 274 888 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3343 0 0
2
5.89796e-315 5.26354e-315
0
13 Logic Switch~
5 342 880 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7923 0 0
2
5.89796e-315 0
0
5 SCOPE
12 476 429 0 1 11
0 3
0
0 0 57584 0
3 TP3
-11 -4 10 4
3 U12
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6174 0 0
2
42835.7 0
0
5 SCOPE
12 473 273 0 1 11
0 4
0
0 0 57584 0
3 TP2
-11 -4 10 4
3 U11
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6692 0 0
2
42835.7 0
0
5 SCOPE
12 169 74 0 1 11
0 5
0
0 0 57584 0
3 TP1
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8790 0 0
2
42835.6 0
0
5 SCOPE
12 98 71 0 1 11
0 6
0
0 0 57584 0
3 CLK
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4595 0 0
2
42835.6 0
0
7 Pulser~
4 563 778 0 10 12
0 36 37 10 38 0 0 10 10 3
8
0
0 0 4656 180
0
2 V3
-7 -29 7 -21
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
667 0 0
2
5.89796e-315 0
0
14 Logic Display~
6 618 780 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8743 0 0
2
5.89796e-315 0
0
7 74LS165
97 405 763 0 14 29
0 8 9 8 9 8 9 8 9 13
12 2 10 39 11
0
0 0 15088 0
7 74LS165
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 0 0 0
1 U
8298 0 0
2
5.89796e-315 5.37752e-315
0
7 Ground~
168 483 735 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
313 0 0
2
5.89796e-315 5.3568e-315
0
7 Pulser~
4 41 94 0 10 12
0 40 41 6 42 0 0 10 10 3
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7548 0 0
2
5.89796e-315 0
0
9 2-In AND~
219 590 536 0 3 22
0 17 16 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8973 0 0
2
5.89796e-315 5.30499e-315
0
7 Ground~
168 167 461 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9712 0 0
2
42835.6 0
0
7 74LS290
153 376 481 0 10 21
0 2 2 14 15 20 18 20 14 3
21
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
2 U7
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
4518 0 0
2
42835.6 1
0
7 74LS290
153 219 482 0 10 21
0 2 2 14 15 19 6 19 16 17
18
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
5596 0 0
2
42835.6 2
0
12 Hex Display~
7 584 453 0 18 19
10 17 16 19 18 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP6
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
692 0 0
2
42835.6 3
0
12 Hex Display~
7 523 454 0 16 19
10 3 14 20 21 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6258 0 0
2
42835.6 4
0
7 Ground~
168 321 447 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5578 0 0
2
42835.6 5
0
9 2-In AND~
219 579 339 0 3 22
0 24 23 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8709 0 0
2
42835.6 6
0
12 Hex Display~
7 573 267 0 18 19
10 24 23 29 25 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9131 0 0
2
42835.6 7
0
12 Hex Display~
7 517 267 0 16 19
10 28 4 27 26 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3645 0 0
2
42835.6 8
0
7 Ground~
168 167 253 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7613 0 0
2
42835.6 9
0
7 Ground~
168 324 241 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9467 0 0
2
42835.6 10
0
7 74LS290
153 369 291 0 10 21
0 2 2 4 22 25 28 26 27 4
28
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
3932 0 0
2
42835.6 11
0
7 74LS290
153 225 289 0 10 21
0 2 2 4 22 6 24 25 29 23
24
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 1 0 0 0
1 U
5288 0 0
2
42835.6 12
0
12 Hex Display~
7 218 51 0 16 19
10 5 30 31 32 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4934 0 0
2
5.89796e-315 5.34643e-315
0
12 Hex Display~
7 262 51 0 18 19
10 7 33 34 35 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5987 0 0
2
5.89796e-315 5.3568e-315
0
7 74LS293
154 346 143 0 8 17
0 7 5 35 5 32 31 30 5
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U2
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
7737 0 0
2
42835.6 13
0
7 74LS293
154 221 143 0 8 17
0 7 5 6 7 35 34 33 7
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U1
-6 15 8 23
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
4200 0 0
2
42835.6 14
0
102
-102335 1 3 0 0 8320 0 0 5 53 0 3
440 439
440 441
476 441
1 -102334 4 0 0 8192 0 6 0 0 77 4
473 285
453 285
453 257
430 257
0 1 5 0 0 4096 0 0 7 92 0 4
227 79
188 79
188 86
169 86
1 0 6 0 0 4096 0 8 0 0 21 2
98 83
98 85
0 0 7 0 0 8192 0 0 0 96 91 3
271 85
279 85
279 113
0 1 8 0 0 8320 0 0 3 10 0 4
368 736
325 736
325 888
286 888
1 0 9 0 0 4224 0 4 0 0 13 3
354 880
354 799
365 799
0 7 8 0 0 0 0 0 11 9 0 3
367 772
367 790
373 790
0 5 8 0 0 0 0 0 11 10 0 3
367 754
367 772
373 772
1 3 8 0 0 0 0 11 11 0 0 4
373 736
367 736
367 754
373 754
2 0 9 0 0 0 0 11 0 0 12 3
373 745
364 745
364 763
4 0 9 0 0 0 0 11 0 0 13 3
373 763
364 763
364 784
8 6 9 0 0 0 0 11 11 0 0 4
373 799
364 799
364 781
373 781
11 1 2 0 0 4096 0 11 12 0 0 4
443 745
466 745
466 729
483 729
3 12 10 0 0 8320 0 9 11 0 0 5
539 785
539 786
445 786
445 754
437 754
14 1 11 0 0 8320 0 11 10 0 0 6
437 799
437 812
557 812
557 813
618 813
618 798
10 1 12 0 0 12432 0 11 2 0 0 6
443 736
444 736
444 698
534 698
534 679
522 679
1 9 13 0 0 8320 0 1 11 0 0 5
529 633
529 649
448 649
448 727
437 727
0 6 6 0 0 4224 0 0 17 20 0 3
100 308
100 509
181 509
0 5 6 0 0 0 0 0 27 21 0 4
100 151
100 308
187 308
187 307
3 3 6 0 0 0 0 13 31 0 0 4
65 85
100 85
100 152
183 152
0 -102334 14 0 0 4096 0 0 0 28 54 2
339 430
282 430
-2659785 0 15 0 0 4096 0 0 0 54 27 3
282 485
327 485
327 479
2 -102270 16 0 0 8320 0 14 0 0 43 3
566 545
559 545
559 505
-102271 1 17 0 0 8192 0 0 14 43 0 3
564 505
566 505
566 527
3 -2659785 15 0 0 0 0 14 0 0 43 3
611 536
618 536
618 505
4 4 15 0 0 12416 0 17 16 0 0 6
187 482
178 482
178 419
327 419
327 481
344 481
3 3 14 0 0 12416 0 17 16 0 0 6
187 473
183 473
183 425
339 425
339 472
344 472
4 -102268 18 0 0 4096 0 18 0 0 43 2
575 477
575 505
1 0 2 0 0 0 0 15 0 0 31 2
167 455
167 455
1 0 2 0 0 0 0 17 0 0 0 2
187 455
164 455
2 1 2 0 0 0 0 17 17 0 0 2
187 464
187 455
5 7 19 0 0 12416 0 17 17 0 0 5
181 500
173 500
173 433
251 433
251 455
7 5 20 0 0 8320 0 16 16 0 0 5
408 454
408 435
334 435
334 499
338 499
1 2 2 0 0 0 0 16 16 0 0 2
344 454
344 463
1 -102271 17 0 0 4096 0 18 0 0 43 2
593 477
593 505
2 -102270 16 0 0 0 0 18 0 0 43 2
587 477
587 505
3 -102269 19 0 0 0 0 18 0 0 43 2
581 477
581 505
1 -102335 3 0 0 128 0 19 0 0 43 2
532 478
532 505
2 -102334 14 0 0 0 0 19 0 0 43 2
526 478
526 505
3 -102333 20 0 0 0 0 19 0 0 43 2
520 478
520 505
4 -102332 21 0 0 4224 0 19 0 0 43 2
514 478
514 505
-407671614 0 1 0 0 4256 0 0 0 0 0 2
477 505
655 505
10 -102332 21 0 0 0 0 16 0 0 53 4
408 508
425 508
425 504
440 504
7 -102333 20 0 0 0 0 16 0 0 53 4
408 454
425 454
425 450
440 450
8 -102334 14 0 0 0 0 16 0 0 53 4
408 472
425 472
425 468
440 468
9 -102335 3 0 0 0 0 16 0 0 53 4
408 490
425 490
425 486
440 486
6 -102268 18 0 0 4224 0 16 0 0 54 4
338 508
303 508
303 519
282 519
10 -102268 18 0 0 0 0 17 0 0 54 2
251 509
282 509
7 -102269 19 0 0 0 0 17 0 0 54 2
251 455
282 455
8 -102270 16 0 0 0 0 17 0 0 54 2
251 473
282 473
9 -102271 17 0 0 4224 0 17 0 0 54 2
251 491
282 491
-407671614 0 1 0 0 32 0 0 0 0 0 2
440 419
440 561
-407671614 0 1 0 0 32 0 0 0 0 0 2
282 413
282 559
1 1 2 0 0 0 0 20 16 0 0 3
321 441
344 441
344 454
0 -2716233 22 0 0 4096 0 0 0 60 82 2
306 290
285 290
3 -2716233 22 0 0 8192 0 21 0 0 72 3
600 339
607 339
607 314
2 -102270 23 0 0 8320 0 21 0 0 72 3
555 348
545 348
545 314
1 -102271 24 0 0 8192 0 21 0 0 72 3
555 330
550 330
550 314
4 4 22 0 0 12416 0 27 26 0 0 6
193 289
183 289
183 226
306 226
306 291
337 291
0 -102334 4 0 0 0 0 0 0 62 82 2
313 250
285 250
3 3 4 0 0 12416 0 26 27 0 0 6
337 282
313 282
313 222
188 222
188 280
193 280
5 -102268 25 0 0 4224 0 26 0 0 82 2
331 309
285 309
4 -102332 26 0 0 4096 0 23 0 0 72 2
508 291
508 314
3 -102333 27 0 0 4096 0 23 0 0 72 2
514 291
514 314
2 -102334 4 0 0 0 0 23 0 0 72 2
520 291
520 314
1 -102335 28 0 0 4096 0 23 0 0 72 2
526 291
526 314
4 -102268 25 0 0 0 0 22 0 0 72 2
564 291
564 314
3 -102269 29 0 0 4096 0 22 0 0 72 2
570 291
570 314
2 -102270 23 0 0 0 0 22 0 0 72 2
576 291
576 314
1 -102271 24 0 0 4096 0 22 0 0 72 2
582 291
582 314
-6369869 0 1 0 0 32 0 0 0 0 0 2
479 314
629 314
10 -102335 28 0 0 4096 0 26 0 0 77 2
401 318
430 318
9 -102334 4 0 0 0 0 26 0 0 77 2
401 300
430 300
8 -102333 27 0 0 4224 0 26 0 0 77 2
401 282
430 282
7 -102332 26 0 0 4224 0 26 0 0 77 2
401 264
430 264
-6369869 0 1 0 0 32 0 0 0 0 0 2
430 234
430 347
10 -102271 24 0 0 4096 0 27 0 0 82 2
257 316
285 316
9 -102270 23 0 0 0 0 27 0 0 82 2
257 298
285 298
8 -102269 29 0 0 4224 0 27 0 0 82 2
257 280
285 280
7 -102268 25 0 0 0 0 27 0 0 82 2
257 262
285 262
-6369869 0 1 0 0 32 0 0 0 0 0 2
285 235
285 348
10 6 28 0 0 8320 0 26 26 0 0 4
401 318
401 330
331 330
331 318
10 6 24 0 0 8320 0 27 27 0 0 4
257 316
257 330
187 330
187 316
1 2 2 0 0 0 0 26 26 0 0 2
337 264
337 273
1 1 2 0 0 8320 0 25 26 0 0 3
324 235
337 235
337 264
1 2 2 0 0 0 0 27 27 0 0 2
193 262
193 271
1 1 2 0 0 0 0 24 27 0 0 3
167 247
193 247
193 262
0 0 5 0 0 0 0 0 0 92 90 3
317 80
291 80
291 109
2 2 5 0 0 12416 0 30 31 0 0 6
314 143
307 143
307 109
183 109
183 143
189 143
1 1 7 0 0 8320 0 31 30 0 0 4
189 134
189 113
314 113
314 134
1 0 5 0 0 0 0 28 0 0 101 7
227 75
227 80
317 80
317 84
394 84
394 161
386 161
2 7 30 0 0 8320 0 28 30 0 0 5
221 75
221 89
390 89
390 152
378 152
6 3 31 0 0 12416 0 30 28 0 0 5
378 143
384 143
384 93
215 93
215 75
5 4 32 0 0 8320 0 30 28 0 0 4
378 134
378 99
209 99
209 75
1 8 7 0 0 128 0 29 31 0 0 3
271 75
271 161
253 161
7 2 33 0 0 8320 0 31 29 0 0 3
253 152
265 152
265 75
3 6 34 0 0 4224 0 29 31 0 0 3
259 75
259 143
253 143
5 4 35 0 0 4224 0 31 29 0 0 2
253 134
253 75
5 3 35 0 0 0 0 31 30 0 0 4
253 134
284 134
284 152
308 152
8 4 5 0 0 0 0 30 30 0 0 5
378 161
387 161
387 179
308 179
308 161
8 4 7 0 0 0 0 31 31 0 0 4
253 161
253 178
183 178
183 161
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 145
-2 610 450 677
15 623 432 675
145 Transforma a informa��o de paralelo para serie.

No circuito abaixo ele alterna entre 1 e 0, at� para 
de acordo com o bit da entrada serial.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
