CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
200 40 30 150 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499450 0.500000
344 176 1846 629
110100498 256
0
6 Title:
5 Name:
0
0
0
19
6 74LS85
106 882 126 0 14 29
0 16 15 5 14 2 2 2 11 20
21 22 41 23 42
0
0 0 5088 0
6 74LS85
-21 -52 21 -44
2 U2
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
331 0 0
2
42847.7 7
0
6 74LS85
106 882 252 0 14 29
0 13 12 4 3 2 2 2 11 38
39 40 20 21 22
0
0 0 5088 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
9604 0 0
2
42847.7 6
0
6 74LS74
17 1089 333 0 12 25
0 23 11 11 10 31 32 33 34 24
35 36 37
0
0 0 4832 0
6 74LS74
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 0 0 0 0
1 U
7518 0 0
2
42847.7 5
0
14 Logic Display~
6 1161 288 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
4 Is11
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4832 0 0
2
42847.7 4
0
2 +V
167 783 63 0 1 3
0 11
0
0 0 53600 0
2 5V
-8 -22 6 -14
3 VCC
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6798 0 0
2
42847.7 3
0
7 Ground~
168 819 603 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3336 0 0
2
42847.7 2
0
6 74LS85
106 882 540 0 14 29
0 13 12 4 3 11 2 2 2 27
28 29 17 18 19
0
0 0 5088 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
8370 0 0
2
42847.7 1
0
6 74LS85
106 882 414 0 14 29
0 16 15 5 14 2 2 2 11 17
18 19 10 25 26
0
0 0 5088 0
6 74LS85
-21 -52 21 -44
2 U6
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3910 0 0
2
42847.7 0
0
13 Logic Switch~
5 225 342 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 Clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
316 0 0
2
42847.7 0
0
13 Logic Switch~
5 234 234 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
7 MasterR
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
536 0 0
2
42847.6 0
0
5 7415~
219 333 324 0 4 22
0 5 4 3 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
4460 0 0
2
42847.7 1
0
8 2-In OR~
219 378 333 0 3 22
0 7 6 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3260 0 0
2
42847.7 0
0
12 Hex Display~
7 540 441 0 16 19
10 14 5 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
7 MaisSIG
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5156 0 0
2
42847.6 2
0
12 Hex Display~
7 612 441 0 16 19
10 3 4 12 13 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
7 MenoSIG
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3133 0 0
2
42847.6 1
0
7 Ground~
168 477 486 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5523 0 0
2
42847.6 0
0
7 Ground~
168 441 324 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3746 0 0
2
42847.6 0
0
7 Ground~
168 522 243 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5668 0 0
2
42847.6 0
0
7 74LS290
153 612 225 0 10 21
0 2 2 9 9 13 14 16 15 5
14
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
7 MaisSIG
-24 -52 25 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 0 0 0 0
1 U
5368 0 0
2
42847.6 0
0
7 74LS290
153 495 315 0 10 21
0 2 2 9 9 8 3 13 12 4
3
0
0 0 4848 0
7 74LS290
-24 -51 25 -43
7 MenoSIG
-24 -52 25 -44
0
15 DVCC=14;DGND=7;
94 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 1 3 12 13 10 11 8 4 5
9 1 3 12 13 10 11 8 4 5
9 0
65 0 0 0 0 0 0 0
1 U
8293 0 0
2
42847.6 0
0
83
12 4 10 0 0 16 0 8 3 0 0 4
914 432
1025 432
1025 324
1051 324
2 0 11 0 0 16 0 3 0 0 44 2
1057 306
783 306
3 0 11 0 0 16 0 3 0 0 44 2
1051 315
783 315
8 0 2 0 0 16 0 7 0 0 43 2
850 576
819 576
7 0 2 0 0 16 0 7 0 0 43 2
850 567
819 567
5 0 11 0 0 16 0 7 0 0 44 2
850 549
783 549
6 0 2 0 0 16 0 7 0 0 43 2
850 558
819 558
5 0 2 0 0 16 0 8 0 0 43 2
850 423
819 423
6 0 2 0 0 16 0 8 0 0 43 2
850 432
819 432
7 0 2 0 0 16 0 8 0 0 43 2
850 441
819 441
8 0 11 0 0 16 0 8 0 0 44 2
850 450
783 450
4 -656179328 3 0 0 16 0 7 0 0 42 2
850 540
743 540
3 -656179327 4 0 0 16 0 7 0 0 42 2
850 531
743 531
2 -656179326 12 0 0 16 0 7 0 0 42 2
850 522
743 522
1 -656179325 13 0 0 16 0 7 0 0 42 2
850 513
743 513
4 -656179324 14 0 0 16 0 8 0 0 42 2
850 414
743 414
3 -656179323 5 0 0 16 0 8 0 0 42 2
850 405
743 405
2 -656179322 15 0 0 16 0 8 0 0 42 2
850 396
743 396
1 -656179321 16 0 0 16 0 8 0 0 42 2
850 387
743 387
9 12 17 0 0 16 0 8 7 0 0 4
914 387
945 387
945 558
914 558
13 10 18 0 0 16 0 7 8 0 0 4
914 567
936 567
936 396
914 396
14 11 19 0 0 16 0 7 8 0 0 4
914 576
928 576
928 405
914 405
3 -656179327 4 0 0 16 0 2 0 0 42 2
850 243
743 243
2 -656179326 12 0 0 16 0 2 0 0 42 2
850 234
743 234
1 -656179325 13 0 0 16 0 2 0 0 42 2
850 225
743 225
3 -656179323 5 0 0 16 0 1 0 0 42 2
850 117
743 117
2 -656179322 15 0 0 16 0 1 0 0 42 2
850 108
743 108
1 -656179321 16 0 0 16 0 1 0 0 42 2
850 99
743 99
5 0 2 0 0 16 0 2 0 0 43 2
850 261
819 261
6 0 2 0 0 16 0 2 0 0 43 2
850 270
819 270
7 0 2 0 0 16 0 2 0 0 43 2
850 279
819 279
8 0 11 0 0 16 0 2 0 0 44 2
850 288
783 288
8 0 11 0 0 16 0 1 0 0 44 2
850 162
783 162
7 0 2 0 0 16 0 1 0 0 43 2
850 153
819 153
6 0 2 0 0 16 0 1 0 0 43 2
850 144
819 144
5 0 2 0 0 16 0 1 0 0 43 2
850 135
819 135
4 -656179328 3 0 0 16 0 2 0 0 42 2
850 252
743 252
4 -656179324 14 0 0 16 0 1 0 0 42 2
850 126
743 126
9 12 20 0 0 16 0 1 2 0 0 4
914 99
945 99
945 270
914 270
13 10 21 0 0 16 0 2 1 0 0 4
914 279
936 279
936 108
914 108
14 11 22 0 0 16 0 2 1 0 0 4
914 288
928 288
928 117
914 117
-594359836 0 1 0 0 48 0 0 0 0 0 2
743 54
743 615
1 0 2 0 0 16 0 6 0 0 0 2
819 597
819 62
1 0 11 0 0 16 0 5 0 0 0 2
783 72
783 612
1 13 23 0 0 16 0 3 1 0 0 4
1057 297
1026 297
1026 153
914 153
9 1 24 0 0 16 0 3 4 0 0 2
1121 306
1161 306
3 -656179328 3 0 0 4096 0 11 0 0 50 2
309 333
261 333
2 -656179327 4 0 0 4096 0 11 0 0 50 2
309 324
261 324
1 -656179323 5 0 0 4096 0 11 0 0 50 2
309 315
261 315
-594359836 0 1 0 0 4128 0 0 0 0 0 2
261 282
261 337
1 2 6 0 0 4224 0 9 12 0 0 2
237 342
365 342
1 4 7 0 0 4224 0 12 11 0 0 2
365 324
354 324
3 5 8 0 0 4224 0 12 19 0 0 2
411 333
457 333
4 0 9 0 0 4096 0 19 0 0 55 3
463 315
451 315
451 306
3 0 9 0 0 8192 0 19 0 0 57 3
463 306
451 306
451 234
4 0 9 0 0 4224 0 18 0 0 57 2
580 225
451 225
1 3 9 0 0 4224 0 10 18 0 0 4
246 234
451 234
451 216
580 216
0 3 9 0 0 0 0 0 19 0 0 2
463 306
463 306
4 0 2 0 0 0 0 13 0 0 60 2
531 465
531 480
3 1 2 0 0 8192 0 13 15 0 0 3
537 465
537 480
477 480
2 -656179323 5 0 0 0 0 13 0 0 67 2
543 465
543 505
1 -656179324 14 0 0 0 0 13 0 0 67 2
549 465
549 505
4 -656179325 13 0 0 0 0 14 0 0 67 2
603 465
603 505
3 -656179326 12 0 0 0 0 14 0 0 67 2
609 465
609 505
2 -656179327 4 0 0 0 0 14 0 0 67 2
615 465
615 505
1 -656179328 3 0 0 0 0 14 0 0 67 2
621 465
621 505
-594359836 0 1 0 0 4128 0 0 0 0 0 2
441 505
679 505
1 0 2 0 0 0 0 19 0 0 69 3
463 288
441 288
441 297
1 2 2 0 0 0 0 16 19 0 0 3
441 318
441 297
463 297
2 0 2 0 0 0 0 18 0 0 71 2
580 207
522 207
1 1 2 0 0 0 0 17 18 0 0 3
522 237
522 198
580 198
0 5 13 0 0 0 0 0 18 79 0 3
540 288
540 243
574 243
0 6 14 0 0 128 0 0 18 78 0 5
657 252
657 271
567 271
567 252
574 252
0 6 3 0 0 0 0 0 19 82 0 5
540 342
540 361
450 361
450 342
457 342
7 -656179321 16 0 0 128 0 18 0 0 83 2
644 198
712 198
8 -656179322 15 0 0 0 0 18 0 0 83 2
644 216
712 216
9 -656179323 5 0 0 128 0 18 0 0 83 2
644 234
712 234
10 -656179324 14 0 0 0 0 18 0 0 83 2
644 252
712 252
7 -656179325 13 0 0 4224 0 19 0 0 83 2
527 288
712 288
8 -656179326 12 0 0 4224 0 19 0 0 83 2
527 306
712 306
9 -656179327 4 0 0 4224 0 19 0 0 83 2
527 324
712 324
10 -656179328 3 0 0 4224 0 19 0 0 83 2
527 342
712 342
-594359836 0 1 0 0 160 0 0 0 0 0 2
712 144
712 386
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
