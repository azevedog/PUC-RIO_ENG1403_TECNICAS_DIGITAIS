CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 130 7 110 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 27 432 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89801e-315 0
0
9 Inverter~
13 765 738 0 2 22
0 4 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
391 0 0
2
42878.4 0
0
12 Hex Display~
7 819 801 0 16 19
10 8 7 6 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
42878.4 0
0
7 Ground~
168 639 918 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3421 0 0
2
42878.4 0
0
7 74LS157
122 702 855 0 14 29
0 3 12 2 11 2 10 2 9 2
2 8 7 6 5
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
8157 0 0
2
42878.4 0
0
7 Ground~
168 648 765 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5572 0 0
2
42878.4 0
0
2 +V
167 630 657 0 1 3
0 13
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
42878.4 0
0
5 4023~
219 477 747 0 4 22
0 9 10 12 14
0
0 0 624 0
4 4023
-14 -28 14 -20
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 4 0
1 U
7361 0 0
2
42878.4 0
0
2 +V
167 288 621 0 1 3
0 16
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
42878.4 0
0
7 Ground~
168 315 729 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
972 0 0
2
42878.4 0
0
7 74LS191
135 396 675 0 14 29
0 2 15 14 2 2 2 38 16 39
40 9 10 11 12
0
0 0 4848 0
7 74LS191
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
3472 0 0
2
42878.4 0
0
12 Hex Display~
7 594 648 0 16 19
10 12 11 10 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9998 0 0
2
5.89801e-315 0
0
5 7415~
219 90 486 0 4 22
0 22 21 36 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
3536 0 0
2
5.89801e-315 0
0
2 +V
167 153 603 0 1 3
0 13
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4597 0 0
2
5.89801e-315 5.26354e-315
0
9 Inverter~
13 540 387 0 2 22
0 25 24
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U6B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3835 0 0
2
5.89801e-315 0
0
2 +V
167 459 396 0 1 3
0 28
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.89801e-315 0
0
7 Ground~
168 486 522 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.89801e-315 0
0
7 74LS190
134 549 459 0 14 29
0 2 23 24 2 2 2 2 2 41
42 43 25 26 27
0
0 0 4848 0
7 74LS190
-24 -51 25 -43
2 U7
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9323 0 0
2
5.89801e-315 0
0
2 +V
167 117 414 0 1 3
0 32
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
5.89801e-315 0
0
9 Inverter~
13 207 423 0 2 22
0 23 33
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U6A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3108 0 0
2
5.89801e-315 0
0
7 74LS190
134 207 495 0 14 29
0 2 15 33 2 2 2 2 32 44
45 46 23 35 34
0
0 0 4848 0
7 74LS190
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4299 0 0
2
5.89801e-315 5.30499e-315
0
7 Ground~
168 144 558 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
5.89801e-315 5.26354e-315
0
6 74LS85
106 702 711 0 14 29
0 9 10 11 12 13 2 13 13 47
48 49 50 4 51
0
0 0 13296 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 79693500
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
5.89801e-315 0
0
7 Ground~
168 729 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
5.89801e-315 0
0
7 Ground~
168 225 374 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
5.89801e-315 0
0
7 74LS153
119 630 243 0 14 29
0 17 29 19 20 26 27 52 53 54
55 2 56 36 57
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
7100 0 0
2
5.89801e-315 0
0
2 +V
167 252 252 0 1 3
0 37
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3820 0 0
2
5.89801e-315 0
0
7 74LS155
120 333 378 0 14 29
0 58 2 35 34 59 60 29 30 31
61 62 63 64 65
0
0 0 4848 0
7 74LS155
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 13 14 15 4 5 6
7 12 11 10 9 1 2 3 13 14
15 4 5 6 7 12 11 10 9 0
65 0 0 512 1 0 0 0
1 U
7678 0 0
2
5.89801e-315 0
0
7 Pulser~
4 29 486 0 10 12
0 66 67 21 68 0 0 10 10 11
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
961 0 0
2
5.89801e-315 0
0
11 4x4 Switch~
193 477 229 0 11 17
0 20 19 29 17 37 29 30 31 0
9 30
0
0 0 4720 512
0
3 SW1
-23 -42 -2 -34
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
2 SW
3178 0 0
2
5.89801e-315 0
0
81
2 1 3 0 0 12416 0 2 5 0 0 6
786 738
801 738
801 759
666 759
666 819
670 819
13 1 4 0 0 4224 0 23 2 0 0 2
734 738
750 738
4 14 5 0 0 8320 0 3 5 0 0 3
810 825
810 891
734 891
3 13 6 0 0 8320 0 3 5 0 0 3
816 825
816 873
734 873
2 12 7 0 0 8320 0 3 5 0 0 3
822 825
822 855
734 855
1 11 8 0 0 8320 0 3 5 0 0 3
828 825
828 837
734 837
3 0 2 0 0 4096 0 5 0 0 12 2
670 837
639 837
5 0 2 0 0 0 0 5 0 0 12 2
670 855
639 855
7 0 2 0 0 0 0 5 0 0 12 2
670 873
639 873
9 0 2 0 0 0 0 5 0 0 12 2
670 891
639 891
10 0 2 0 0 0 0 5 0 0 12 2
664 900
639 900
1 0 2 0 0 4224 0 4 0 0 0 2
639 912
639 801
0 8 9 0 0 4224 0 0 5 26 0 3
586 684
586 882
670 882
0 6 10 0 0 4224 0 0 5 25 0 3
591 693
591 864
670 864
0 4 11 0 0 4096 0 0 5 24 0 3
597 702
597 846
670 846
0 2 12 0 0 4096 0 0 5 23 0 3
604 711
604 828
670 828
6 0 2 0 0 0 0 23 0 0 21 2
670 729
648 729
8 0 13 0 0 4096 0 23 0 0 22 2
670 747
630 747
7 0 13 0 0 0 0 23 0 0 22 2
670 738
630 738
5 0 13 0 0 0 0 23 0 0 22 2
670 720
630 720
1 0 2 0 0 0 0 6 0 0 0 2
648 759
648 667
1 0 13 0 0 4224 0 7 0 0 0 2
630 666
630 756
0 4 12 0 0 0 0 0 23 34 0 2
603 711
670 711
0 3 11 0 0 0 0 0 23 33 0 2
597 702
670 702
0 2 10 0 0 0 0 0 23 32 0 2
591 693
670 693
0 1 9 0 0 0 0 0 23 31 0 2
585 684
670 684
3 0 12 0 0 0 0 8 0 0 34 3
453 756
432 756
432 711
2 0 10 0 0 0 0 8 0 0 32 3
453 747
442 747
442 693
1 0 9 0 0 0 0 8 0 0 31 2
453 738
453 684
4 3 14 0 0 12416 0 8 11 0 0 6
504 747
505 747
505 774
342 774
342 666
358 666
11 4 9 0 0 128 0 11 12 0 0 3
428 684
585 684
585 672
12 3 10 0 0 128 0 11 12 0 0 3
428 693
591 693
591 672
13 2 11 0 0 4224 0 11 12 0 0 3
428 702
597 702
597 672
14 1 12 0 0 4224 0 11 12 0 0 3
428 711
603 711
603 672
0 2 15 0 0 8320 0 0 11 50 0 3
132 486
132 657
364 657
1 0 2 0 0 0 0 11 0 0 43 2
358 648
315 648
4 0 2 0 0 0 0 11 0 0 43 2
364 675
315 675
5 0 2 0 0 0 0 11 0 0 43 2
364 684
315 684
6 0 2 0 0 0 0 11 0 0 43 2
364 693
315 693
0 0 2 0 0 0 0 0 0 0 43 2
371 701
315 701
8 0 16 0 0 4096 0 11 0 0 42 2
364 711
288 711
1 0 16 0 0 4224 0 9 0 0 0 2
288 630
288 729
1 0 2 0 0 0 0 10 0 0 0 2
315 723
315 630
1 4 17 0 0 12416 0 26 30 0 0 6
598 207
592 207
592 198
525 198
525 251
510 251
2 3 29 0 0 12416 18 26 30 0 0 4
598 216
559 216
559 236
510 236
2 3 19 0 0 4224 0 30 26 0 0 4
510 222
578 222
578 225
598 225
4 1 20 0 0 12416 0 26 30 0 0 4
598 234
585 234
585 207
510 207
3 2 21 0 0 4224 0 29 13 0 0 4
53 477
62 477
62 486
66 486
1 1 22 0 0 4224 0 13 1 0 0 3
66 477
66 432
39 432
4 2 15 0 0 0 0 13 21 0 0 4
111 486
132 486
132 477
175 477
0 2 23 0 0 12416 0 0 18 69 0 4
253 513
381 513
381 441
517 441
2 3 24 0 0 8320 0 15 18 0 0 4
525 387
504 387
504 450
511 450
12 1 25 0 0 8320 0 18 15 0 0 6
581 477
591 477
591 397
566 397
566 387
561 387
13 5 26 0 0 8320 0 18 26 0 0 6
581 486
602 486
602 343
566 343
566 243
598 243
14 6 27 0 0 8320 0 18 26 0 0 6
581 495
614 495
614 332
576 332
576 252
598 252
8 0 2 0 0 0 0 18 0 0 63 2
517 495
486 495
7 0 2 0 0 0 0 18 0 0 63 2
517 486
486 486
6 0 2 0 0 0 0 18 0 0 63 2
517 477
486 477
5 0 2 0 0 0 0 18 0 0 63 2
517 468
486 468
4 0 2 0 0 0 0 18 0 0 63 2
517 459
486 459
1 0 2 0 0 0 0 18 0 0 63 2
511 432
486 432
1 0 28 0 0 4224 0 16 0 0 0 2
459 405
459 522
1 0 2 0 0 128 0 17 0 0 0 2
486 516
486 409
7 6 29 0 0 4224 0 28 30 0 0 3
371 351
481 351
481 280
8 7 30 0 0 4224 0 28 30 0 0 3
371 360
466 360
466 280
9 8 31 0 0 8320 0 28 30 0 0 3
371 369
452 369
452 280
8 1 32 0 0 8320 0 21 19 0 0 3
175 531
117 531
117 423
2 3 33 0 0 8320 0 20 21 0 0 4
192 423
157 423
157 486
169 486
12 1 23 0 0 0 0 21 20 0 0 4
239 513
253 513
253 423
228 423
14 4 34 0 0 8320 0 21 28 0 0 4
239 531
288 531
288 387
301 387
13 3 35 0 0 8320 0 21 28 0 0 4
239 522
279 522
279 378
301 378
1 0 2 0 0 0 0 21 0 0 77 2
169 468
144 468
4 0 2 0 0 0 0 21 0 0 77 2
175 495
144 495
7 0 2 0 0 0 0 21 0 0 77 2
175 522
144 522
6 0 2 0 0 0 0 21 0 0 77 2
175 513
144 513
5 0 2 0 0 0 0 21 0 0 77 2
175 504
144 504
1 0 2 0 0 0 0 22 0 0 0 2
144 552
144 445
11 1 2 0 0 0 0 26 24 0 0 5
668 207
692 207
692 135
729 135
729 165
1 2 2 0 0 0 0 25 28 0 0 3
225 368
225 360
295 360
3 13 36 0 0 8320 0 13 26 0 0 7
66 495
66 595
650 595
650 352
718 352
718 225
662 225
5 1 37 0 0 8320 0 30 27 0 0 4
437 280
437 315
252 315
252 261
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
