CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
110 270 30 130 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 281 515 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 Clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
313 0 0
2
42847.8 1
0
13 Logic Switch~
5 281 452 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 MODO
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7548 0 0
2
42847.8 0
0
9 2-In AND~
219 1062 567 0 3 22
0 11 4 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8973 0 0
2
42847.8 0
0
6 74LS85
106 922 362 0 14 29
0 10 9 8 7 2 2 2 6 19
20 21 11 37 38
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U2
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9712 0 0
2
42847.8 6
0
6 74LS85
106 922 488 0 14 29
0 15 14 13 12 6 2 2 2 39
40 41 19 20 21
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4518 0 0
2
42847.8 5
0
2 +V
167 823 299 0 1 3
0 6
0
0 0 53616 0
2 5V
-8 -22 6 -14
3 VCC
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5596 0 0
2
42847.8 4
0
7 Ground~
168 859 839 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
692 0 0
2
42847.8 3
0
6 74LS85
106 922 776 0 14 29
0 15 14 13 12 2 6 2 6 42
43 44 16 17 18
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6258 0 0
2
42847.8 2
0
6 74LS85
106 922 650 0 14 29
0 10 9 8 7 2 2 2 2 16
17 18 45 46 4
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U6
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5578 0 0
2
42847.8 1
0
7 74LS157
122 630 855 0 14 29
0 4 2 2 5 5 5 5 5 2
2 25 24 23 22
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8709 0 0
2
42847.8 3
0
7 74LS157
122 630 738 0 14 29
0 4 2 2 2 2 2 2 5 2
2 29 28 27 26
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9131 0 0
2
42847.8 2
0
2 +V
167 535 686 0 1 3
0 5
0
0 0 53616 0
2 5V
-8 -22 6 -14
4 VCC1
-13 -32 15 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3645 0 0
2
42847.8 1
0
7 Ground~
168 562 920 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7613 0 0
2
42847.8 0
0
7 Ground~
168 333 549 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9467 0 0
2
42847.8 10
0
2 +V
167 315 477 0 1 3
0 34
0
0 0 53616 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3932 0 0
2
42847.8 9
0
7 74LS157
122 378 486 0 14 29
0 36 47 48 49 50 34 35 35 34
2 51 52 33 32
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
5288 0 0
2
42847.8 8
0
7 74LS193
137 517 531 0 14 29
0 33 32 3 2 25 24 23 22 30
31 15 14 13 12
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 0 1 0 0 0
1 U
4934 0 0
2
42847.8 7
0
7 Ground~
168 432 585 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5987 0 0
2
42847.8 6
0
7 Ground~
168 621 603 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7737 0 0
2
42847.8 5
0
7 74LS193
137 715 549 0 14 29
0 30 31 3 2 29 28 27 26 53
54 10 9 8 7
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4200 0 0
2
42847.8 4
0
12 Hex Display~
7 315 603 0 16 19
10 7 8 9 10 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5780 0 0
2
42847.8 3
0
12 Hex Display~
7 369 603 0 18 19
10 12 13 14 15 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6490 0 0
2
42847.8 2
0
119
0 -13423565 3 0 0 4096 0 0 0 30 2 2
469 469
432 469
-2475 0 1 0 0 4144 0 0 0 0 0 2
432 436
432 488
1 0 4 0 0 4096 0 10 0 0 4 2
598 819
585 819
0 1 4 0 0 8320 0 0 11 31 0 5
1009 686
1009 919
585 919
585 702
598 702
8 0 5 0 0 4096 0 10 0 0 83 2
598 882
535 882
6 0 5 0 0 0 0 10 0 0 83 2
598 864
535 864
4 0 5 0 0 0 0 10 0 0 83 2
598 846
535 846
2 0 2 0 0 4096 0 10 0 0 82 2
598 828
562 828
8 0 5 0 0 0 0 11 0 0 83 2
598 765
535 765
6 0 2 0 0 0 0 11 0 0 82 2
598 747
562 747
4 0 2 0 0 0 0 11 0 0 82 2
598 729
562 729
2 0 2 0 0 0 0 11 0 0 82 2
598 711
562 711
10 0 2 0 0 0 0 11 0 0 82 2
592 783
562 783
10 0 2 0 0 0 0 10 0 0 82 2
592 900
562 900
9 0 2 0 0 0 0 10 0 0 82 2
598 891
562 891
7 0 5 0 0 0 0 10 0 0 83 2
598 873
535 873
5 0 5 0 0 0 0 10 0 0 83 2
598 855
535 855
3 0 2 0 0 0 0 10 0 0 82 2
598 837
562 837
9 0 2 0 0 0 0 11 0 0 82 2
598 774
562 774
7 0 2 0 0 0 0 11 0 0 82 2
598 756
562 756
5 0 2 0 0 0 0 11 0 0 82 2
598 738
562 738
3 0 2 0 0 0 0 11 0 0 82 2
598 720
562 720
8 0 6 0 0 4096 0 8 0 0 72 2
890 812
823 812
7 0 2 0 0 0 0 8 0 0 71 2
890 803
859 803
6 0 6 0 0 0 0 8 0 0 72 2
890 794
823 794
8 0 2 0 0 0 0 5 0 0 71 2
890 524
859 524
7 0 2 0 0 0 0 5 0 0 71 2
890 515
859 515
6 0 2 0 0 0 0 5 0 0 71 2
890 506
859 506
5 0 6 0 0 0 0 5 0 0 72 2
890 497
823 497
3 3 3 0 0 12416 0 17 20 0 0 6
479 522
469 522
469 469
667 469
667 540
677 540
14 2 4 0 0 128 0 9 3 0 0 4
954 686
1009 686
1009 576
1038 576
14 -656179324 7 0 0 4096 0 20 0 0 70 2
747 585
783 585
13 -656179323 8 0 0 4096 0 20 0 0 70 2
747 576
783 576
12 -656179322 9 0 0 4096 0 20 0 0 70 2
747 567
783 567
11 -656179321 10 0 0 4096 0 20 0 0 70 2
747 558
783 558
3 -13423565 3 0 0 128 0 3 0 0 37 2
1083 567
1134 567
-2475 0 1 0 0 32 0 0 0 0 0 2
1134 535
1134 587
12 1 11 0 0 8320 0 4 3 0 0 4
954 380
1009 380
1009 558
1038 558
5 0 2 0 0 0 0 8 0 0 71 2
890 785
859 785
8 0 2 0 0 0 0 9 0 0 71 2
890 686
859 686
5 0 2 0 0 0 0 9 0 0 71 2
890 659
859 659
6 0 2 0 0 0 0 9 0 0 71 2
890 668
859 668
7 0 2 0 0 0 0 9 0 0 71 2
890 677
859 677
4 -656179328 12 0 0 4224 0 8 0 0 70 2
890 776
783 776
3 -656179327 13 0 0 4224 0 8 0 0 70 2
890 767
783 767
2 -656179326 14 0 0 4224 0 8 0 0 70 2
890 758
783 758
1 -656179325 15 0 0 4224 0 8 0 0 70 2
890 749
783 749
4 -656179324 7 0 0 4224 0 9 0 0 70 2
890 650
783 650
3 -656179323 8 0 0 4224 0 9 0 0 70 2
890 641
783 641
2 -656179322 9 0 0 4224 0 9 0 0 70 2
890 632
783 632
1 -656179321 10 0 0 4224 0 9 0 0 70 2
890 623
783 623
9 12 16 0 0 8320 0 9 8 0 0 4
954 623
985 623
985 794
954 794
13 10 17 0 0 8320 0 8 9 0 0 4
954 803
976 803
976 632
954 632
14 11 18 0 0 8320 0 8 9 0 0 4
954 812
968 812
968 641
954 641
3 -656179327 13 0 0 0 0 5 0 0 70 2
890 479
783 479
2 -656179326 14 0 0 0 0 5 0 0 70 2
890 470
783 470
1 -656179325 15 0 0 0 0 5 0 0 70 2
890 461
783 461
3 -656179323 8 0 0 0 0 4 0 0 70 2
890 353
783 353
2 -656179322 9 0 0 0 0 4 0 0 70 2
890 344
783 344
1 -656179321 10 0 0 0 0 4 0 0 70 2
890 335
783 335
8 0 6 0 0 0 0 4 0 0 72 2
890 398
823 398
7 0 2 0 0 0 0 4 0 0 71 2
890 389
859 389
6 0 2 0 0 0 0 4 0 0 71 2
890 380
859 380
5 0 2 0 0 0 0 4 0 0 71 2
890 371
859 371
4 -656179328 12 0 0 0 0 5 0 0 70 2
890 488
783 488
4 -656179324 7 0 0 0 0 4 0 0 70 2
890 362
783 362
9 12 19 0 0 8320 0 4 5 0 0 4
954 335
985 335
985 506
954 506
13 10 20 0 0 8320 0 5 4 0 0 4
954 515
976 515
976 344
954 344
14 11 21 0 0 8320 0 5 4 0 0 4
954 524
968 524
968 353
954 353
-160201 0 1 0 0 4256 0 0 0 0 0 2
783 290
783 851
1 0 2 0 0 4224 0 7 0 0 0 2
859 833
859 298
1 0 6 0 0 4224 0 6 0 0 0 2
823 308
823 848
14 -143488 22 0 0 4224 0 10 0 0 81 2
662 891
721 891
13 -143487 23 0 0 4224 0 10 0 0 81 2
662 873
721 873
12 -143486 24 0 0 4224 0 10 0 0 81 2
662 855
721 855
11 -143485 25 0 0 4224 0 10 0 0 81 2
662 837
721 837
14 -143484 26 0 0 4224 0 11 0 0 81 2
662 774
721 774
13 -143483 27 0 0 4224 0 11 0 0 81 2
662 756
721 756
12 -143482 28 0 0 4224 0 11 0 0 81 2
662 738
721 738
11 -143481 29 0 0 4224 0 11 0 0 81 2
662 720
721 720
-144841 0 1 0 0 32 0 0 0 0 0 2
721 683
721 911
1 0 2 0 0 0 0 13 0 0 0 2
562 914
562 684
1 0 5 0 0 4224 0 12 0 0 0 2
535 695
535 919
8 -143484 26 0 0 0 0 20 0 0 88 2
683 585
649 585
7 -143483 27 0 0 0 0 20 0 0 88 2
683 576
649 576
6 -143482 28 0 0 0 0 20 0 0 88 2
683 567
649 567
5 -143481 29 0 0 0 0 20 0 0 88 2
683 558
649 558
-144841 0 1 0 0 32 0 0 0 0 0 2
649 627
649 553
8 -143488 22 0 0 0 0 17 0 0 93 2
485 567
451 567
7 -143487 23 0 0 0 0 17 0 0 93 2
485 558
451 558
6 -143486 24 0 0 0 0 17 0 0 93 2
485 549
451 549
5 -143485 25 0 0 0 0 17 0 0 93 2
485 540
451 540
-144841 0 1 0 0 32 0 0 0 0 0 2
451 611
451 536
1 4 2 0 0 0 0 19 20 0 0 3
621 597
621 549
683 549
4 1 2 0 0 0 0 17 18 0 0 3
485 531
432 531
432 579
4 -656179321 10 0 0 0 0 21 0 0 104 2
306 627
306 674
3 -656179322 9 0 0 0 0 21 0 0 104 2
312 627
312 674
2 -656179323 8 0 0 0 0 21 0 0 104 2
318 627
318 674
1 -656179324 7 0 0 0 0 21 0 0 104 2
324 627
324 674
4 -656179325 15 0 0 0 0 22 0 0 104 2
360 627
360 674
3 -656179326 14 0 0 0 0 22 0 0 104 2
366 627
366 674
2 -656179327 13 0 0 0 0 22 0 0 104 2
372 627
372 674
-656179328 1 12 0 0 0 0 0 22 104 0 2
378 674
378 627
-160201 0 1 0 0 32 0 0 0 0 0 2
405 674
279 674
9 1 30 0 0 4224 0 17 20 0 0 2
555 522
683 522
-160201 0 1 0 0 32 0 0 0 0 0 2
595 631
595 535
10 2 31 0 0 4224 0 17 20 0 0 2
555 531
683 531
14 2 32 0 0 12416 0 16 17 0 0 4
410 522
424 522
424 513
485 513
1 13 33 0 0 4224 0 17 16 0 0 2
485 504
410 504
14 -656179328 12 0 0 0 0 17 0 0 106 2
549 567
595 567
13 -656179327 13 0 0 0 0 17 0 0 106 2
549 558
595 558
12 -656179326 14 0 0 0 0 17 0 0 106 2
549 549
595 549
11 -656179325 15 0 0 0 0 17 0 0 106 2
549 540
595 540
0 9 34 0 0 8320 0 0 16 115 0 3
315 495
315 522
346 522
1 6 34 0 0 0 0 15 16 0 0 3
315 486
315 495
346 495
0 1 35 0 0 8320 0 0 1 117 0 3
325 513
325 515
293 515
7 8 35 0 0 0 0 16 16 0 0 4
346 504
325 504
325 513
346 513
10 1 2 0 0 0 0 16 14 0 0 3
340 531
333 531
333 543
1 1 36 0 0 8320 0 16 2 0 0 3
346 450
346 452
293 452
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
