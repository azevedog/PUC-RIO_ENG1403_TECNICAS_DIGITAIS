CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 90 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
40
2 +V
167 651 196 0 1 3
0 25
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
361 0 0
2
42834.7 0
0
7 Ground~
168 872 207 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3343 0 0
2
5.89796e-315 0
0
12 Hex Display~
7 896 177 0 16 19
10 4 5 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7923 0 0
2
5.89796e-315 0
0
7 Ground~
168 861 265 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6174 0 0
2
5.89796e-315 0
0
12 Hex Display~
7 944 254 0 16 19
10 13 12 11 10 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 Alarm
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6692 0 0
2
5.89796e-315 0
0
12 Hex Display~
7 894 256 0 16 19
10 9 2 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 Temp
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8790 0 0
2
5.89796e-315 0
0
7 Ground~
168 745 481 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4595 0 0
2
5.89796e-315 0
0
7 74LS157
122 793 431 0 14 29
0 8 14 2 7 2 6 2 2 2
2 9 4 5 60
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
3 U14
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
667 0 0
2
5.89796e-315 0
0
7 Ground~
168 745 363 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8743 0 0
2
5.89796e-315 0
0
7 74LS157
122 789 312 0 14 29
0 8 18 2 17 2 16 2 15 2
2 13 12 11 10
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
3 U13
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8298 0 0
2
5.89796e-315 0
0
12 Hex Display~
7 591 367 0 16 19
10 14 61 62 63 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 Temp
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
313 0 0
2
5.89796e-315 0
0
7 Ground~
168 489 627 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7548 0 0
2
42834.7 0
0
6 74LS83
105 566 514 0 14 29
0 20 21 22 23 2 19 19 2 2
15 16 17 18 14
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U11
-11 -61 10 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8973 0 0
2
42834.7 1
0
2 +V
167 348 553 0 1 3
0 24
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9712 0 0
2
42834.7 2
0
7 Ground~
168 358 578 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4518 0 0
2
42834.7 3
0
6 74LS85
106 405 525 0 14 29
0 20 21 22 23 24 2 2 24 64
65 66 67 68 19
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
3 U10
-10 -62 11 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5596 0 0
2
42834.7 4
0
6 74LS93
109 319 91 0 8 17
0 26 26 3 7 27 26 6 7
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U9
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
692 0 0
2
42834.7 6
0
7 Pulser~
4 195 26 0 10 12
0 69 70 3 71 0 0 10 10 2
7
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6258 0 0
2
42834.7 7
0
12 Hex Display~
7 414 53 0 16 19
10 7 6 26 27 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5578 0 0
2
42834.7 8
0
14 Logic Display~
6 773 150 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 ALARM
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8709 0 0
2
5.89796e-315 0
0
6 74LS74
17 704 153 0 12 25
0 72 73 74 75 3 8 25 25 76
77 28 78
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U8
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 1 0 0 0
1 U
9131 0 0
2
5.89796e-315 5.26354e-315
0
7 Ground~
168 495 331 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3645 0 0
2
5.89796e-315 5.32571e-315
0
12 Hex Display~
7 616 282 0 16 19
10 7 6 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 NTanq
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7613 0 0
2
5.89796e-315 5.34643e-315
0
2 +V
167 434 163 0 1 3
0 29
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9467 0 0
2
5.89796e-315 5.3568e-315
0
7 Ground~
168 485 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3932 0 0
2
5.89796e-315 5.36716e-315
0
6 74LS85
106 539 152 0 14 29
0 20 21 22 23 29 2 29 29 79
80 81 82 83 8
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U7
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5288 0 0
2
5.89796e-315 5.37752e-315
0
9 2-In AND~
219 317 299 0 3 22
0 7 6 38
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U6A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4934 0 0
2
5.89796e-315 5.38788e-315
0
8 2-In OR~
219 273 174 0 3 22
0 42 41 39
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5987 0 0
2
5.89796e-315 5.39306e-315
0
7 Ground~
168 345 451 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7737 0 0
2
5.89796e-315 5.39824e-315
0
7 74LS157
122 395 400 0 14 29
0 39 46 50 45 49 44 48 43 47
2 23 22 21 20
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
4200 0 0
2
5.89796e-315 5.40342e-315
0
12 Hex Display~
7 636 367 0 16 19
10 18 17 16 15 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 Decim
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5780 0 0
2
5.89796e-315 5.4086e-315
0
2 +V
167 48 144 0 1 3
0 51
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6490 0 0
2
5.89796e-315 5.41378e-315
0
7 Ground~
168 137 247 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8663 0 0
2
5.89796e-315 5.41896e-315
0
7 74LS157
122 233 340 0 14 29
0 7 55 59 54 58 53 57 52 56
39 50 49 48 47
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
318 0 0
2
5.89796e-315 5.42414e-315
0
7 74LS157
122 234 493 0 14 29
0 38 33 37 32 36 31 35 30 34
40 46 45 44 43
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
348 0 0
2
5.89796e-315 5.42933e-315
0
8 Hex Key~
166 66 287 0 11 12
0 59 58 57 56 0 0 0 0 0
0 48
0
0 0 4656 0
0
5 Temp0
-17 -34 18 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8551 0 0
2
5.89796e-315 5.43192e-315
0
8 Hex Key~
166 65 376 0 11 12
0 55 54 53 52 0 0 0 0 0
1 49
0
0 0 4656 0
0
5 Temp1
-17 -34 18 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7295 0 0
2
5.89796e-315 5.43451e-315
0
8 Hex Key~
166 64 471 0 11 12
0 37 36 35 34 0 0 0 0 0
2 50
0
0 0 4656 0
0
5 Temp2
-17 -34 18 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9900 0 0
2
5.89796e-315 5.4371e-315
0
8 Hex Key~
166 61 555 0 11 12
0 33 32 31 30 0 0 0 0 0
12 67
0
0 0 4656 0
0
5 Temp3
-17 -34 18 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8725 0 0
2
5.89796e-315 5.43969e-315
0
6 74LS85
106 182 130 0 14 29
0 2 2 6 7 2 2 51 2 84
85 86 40 42 41
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
366 0 0
2
5.89796e-315 5.44228e-315
0
124
0 5 3 0 0 4224 0 0 21 64 0 4
279 18
626 18
626 162
672 162
5 3 2 0 0 4096 0 8 8 0 0 2
761 431
761 413
12 1 4 0 0 8320 0 8 3 0 0 5
825 431
846 431
846 214
905 214
905 201
2 13 5 0 0 12416 0 3 8 0 0 5
899 201
899 217
855 217
855 449
825 449
1 0 2 0 0 0 0 2 0 0 6 2
872 201
872 201
4 0 2 0 0 0 0 3 0 0 0 2
887 201
869 201
3 4 2 0 0 0 0 3 3 0 0 2
893 201
887 201
8 9 2 0 0 0 0 8 8 0 0 2
761 458
761 467
7 8 2 0 0 0 0 8 8 0 0 2
761 449
761 458
5 7 2 0 0 0 0 8 8 0 0 2
761 431
761 449
6 2 6 0 0 16384 0 8 23 0 0 6
761 440
722 440
722 443
663 443
663 306
619 306
0 4 7 0 0 8192 0 0 8 77 0 4
623 323
675 323
675 422
761 422
0 0 8 0 0 8192 0 0 0 14 34 4
627 188
627 243
719 243
719 277
14 6 8 0 0 0 0 26 21 0 0 4
571 188
627 188
627 171
672 171
9 0 2 0 0 0 0 8 0 0 35 3
761 467
752 467
752 476
1 0 2 0 0 0 0 4 0 0 17 2
861 259
861 260
4 0 2 0 0 8192 0 6 0 0 0 4
885 280
873 280
873 260
857 260
3 4 2 0 0 0 0 6 6 0 0 2
891 280
885 280
2 3 2 0 0 0 0 6 6 0 0 2
897 280
891 280
11 1 9 0 0 8320 0 8 6 0 0 3
825 413
903 413
903 280
4 14 10 0 0 8320 0 5 10 0 0 3
935 278
935 348
821 348
3 13 11 0 0 8320 0 5 10 0 0 3
941 278
941 330
821 330
2 12 12 0 0 8320 0 5 10 0 0 3
947 278
947 312
821 312
11 1 13 0 0 4224 0 10 5 0 0 3
821 294
953 294
953 278
2 0 14 0 0 16384 0 8 0 0 50 5
761 404
761 407
711 407
711 439
600 439
8 0 15 0 0 8192 0 10 0 0 43 4
757 339
685 339
685 431
627 431
6 0 16 0 0 8192 0 10 0 0 42 4
757 321
695 321
695 419
633 419
4 0 17 0 0 8192 0 10 0 0 41 4
757 303
702 303
702 406
639 406
2 0 18 0 0 8192 0 10 0 0 40 4
757 285
706 285
706 396
645 396
0 10 2 0 0 0 0 0 10 31 0 3
750 348
751 348
751 357
0 9 2 0 0 0 0 0 10 32 0 3
750 329
750 348
757 348
0 7 2 0 0 0 0 0 10 33 0 3
750 312
750 330
757 330
3 5 2 0 0 0 0 10 10 0 0 4
757 294
750 294
750 312
757 312
1 1 8 0 0 8320 0 8 10 0 0 4
761 395
719 395
719 276
757 276
1 10 2 0 0 0 0 7 8 0 0 3
745 475
745 476
755 476
1 10 2 0 0 0 0 9 10 0 0 2
745 357
751 357
8 0 2 0 0 8192 0 13 0 0 49 4
534 541
517 541
517 580
515 580
6 7 19 0 0 4096 0 13 13 0 0 4
534 523
534 567
534 567
534 532
7 6 2 0 0 0 0 16 16 0 0 2
373 552
373 543
1 13 18 0 0 4224 0 31 13 0 0 3
645 391
645 532
598 532
12 2 17 0 0 8320 0 13 31 0 0 3
598 523
639 523
639 391
3 11 16 0 0 4224 0 31 13 0 0 3
633 391
633 514
598 514
10 4 15 0 0 8320 0 13 31 0 0 3
598 505
627 505
627 391
14 6 19 0 0 4224 0 16 13 0 0 3
437 561
534 561
534 523
1 0 20 0 0 8192 0 13 0 0 58 3
534 478
534 446
449 446
0 2 21 0 0 4096 0 0 13 57 0 4
452 428
515 428
515 487
534 487
3 0 22 0 0 8192 0 13 0 0 55 4
534 496
510 496
510 410
457 410
0 4 23 0 0 8192 0 0 13 54 0 4
469 455
504 455
504 505
534 505
5 0 2 0 0 8192 0 13 0 0 51 3
534 514
515 514
515 598
1 14 14 0 0 4224 0 11 13 0 0 3
600 391
600 559
598 559
1 9 2 0 0 0 0 12 13 0 0 5
489 621
489 598
515 598
515 559
534 559
14 0 20 0 0 0 0 30 0 0 58 3
427 436
427 446
438 446
13 0 21 0 0 0 0 30 0 0 57 3
427 418
427 428
443 428
0 4 23 0 0 8192 0 0 16 56 0 5
469 380
469 458
356 458
356 525
373 525
0 3 22 0 0 8192 0 0 16 80 0 5
457 409
457 464
362 464
362 516
373 516
4 11 23 0 0 8320 0 26 30 0 0 4
507 152
469 152
469 382
427 382
2 2 21 0 0 24704 0 16 26 0 0 8
373 507
369 507
369 472
443 472
443 428
453 428
453 134
507 134
1 1 20 0 0 8320 0 26 16 0 0 7
507 125
449 125
449 446
438 446
438 477
373 477
373 498
0 1 24 0 0 8192 0 0 14 61 0 3
364 560
364 562
348 562
6 1 2 0 0 0 0 16 15 0 0 3
373 543
358 543
358 572
5 8 24 0 0 8320 0 16 16 0 0 4
373 534
364 534
364 561
373 561
8 1 25 0 0 4224 0 21 1 0 0 4
666 189
666 206
651 206
651 205
7 8 25 0 0 0 0 21 21 0 0 2
666 180
666 189
3 3 3 0 0 128 0 17 18 0 0 4
281 100
279 100
279 17
219 17
4 0 7 0 0 16512 0 40 0 0 95 5
150 130
118 130
118 61
256 61
256 264
0 0 6 0 0 0 0 0 0 71 94 4
398 100
398 219
289 219
289 273
0 0 7 0 0 0 0 0 0 72 95 4
378 109
378 232
324 232
324 264
0 1 26 0 0 8320 0 0 17 70 0 4
362 92
362 54
287 54
287 82
5 4 27 0 0 4224 0 17 19 0 0 3
351 82
405 82
405 77
3 6 26 0 0 0 0 19 17 0 0 5
411 77
411 92
362 92
362 91
351 91
7 2 6 0 0 0 0 17 19 0 0 3
351 100
417 100
417 77
1 8 7 0 0 0 0 19 17 0 0 3
423 77
423 109
351 109
2 1 26 0 0 0 0 17 17 0 0 2
287 91
287 82
8 4 7 0 0 0 0 17 17 0 0 4
351 109
351 122
281 122
281 109
11 1 28 0 0 4224 0 21 20 0 0 3
736 171
773 171
773 168
2 2 6 0 0 4224 0 23 27 0 0 4
619 306
394 306
394 290
335 290
0 1 7 0 0 0 0 0 23 95 0 5
347 307
469 307
469 323
625 323
625 306
4 1 2 0 0 4224 0 23 22 0 0 3
607 306
495 306
495 325
3 4 2 0 0 0 0 23 23 0 0 4
613 306
526 306
526 306
607 306
3 12 22 0 0 8320 0 26 30 0 0 5
507 143
457 143
457 410
427 410
427 400
7 1 29 0 0 4224 0 26 24 0 0 3
507 179
434 179
434 172
8 7 29 0 0 0 0 26 26 0 0 2
507 188
507 179
5 7 29 0 0 0 0 26 26 0 0 4
507 161
501 161
501 179
507 179
6 1 2 0 0 0 0 26 25 0 0 3
507 170
485 170
485 197
4 8 30 0 0 8320 0 39 35 0 0 5
52 579
52 590
165 590
165 520
202 520
6 3 31 0 0 12416 0 35 39 0 0 5
202 502
173 502
173 586
58 586
58 579
2 4 32 0 0 8320 0 39 35 0 0 5
64 579
64 583
179 583
179 484
202 484
2 1 33 0 0 12416 0 35 39 0 0 4
202 466
184 466
184 579
70 579
4 9 34 0 0 16512 0 38 35 0 0 5
55 495
55 517
82 517
82 529
202 529
7 3 35 0 0 4224 0 35 38 0 0 3
202 511
61 511
61 495
2 5 36 0 0 16512 0 38 35 0 0 5
67 495
67 499
88 499
88 493
202 493
3 1 37 0 0 4224 0 35 38 0 0 4
202 475
82 475
82 495
73 495
3 1 38 0 0 8320 0 27 35 0 0 6
290 299
269 299
269 423
195 423
195 457
202 457
3 2 6 0 0 0 0 40 27 0 0 7
150 121
106 121
106 70
239 70
239 273
335 273
335 290
1 1 7 0 0 0 0 34 27 0 0 5
201 304
201 264
347 264
347 308
335 308
3 1 39 0 0 8320 0 28 30 0 0 4
306 174
361 174
361 364
363 364
12 10 40 0 0 16512 0 40 35 0 0 6
214 148
227 148
227 233
191 233
191 538
196 538
3 10 39 0 0 0 0 28 34 0 0 5
306 174
306 201
145 201
145 385
195 385
14 2 41 0 0 12416 0 40 28 0 0 4
214 166
221 166
221 183
260 183
13 1 42 0 0 4224 0 40 28 0 0 4
214 157
253 157
253 165
260 165
10 1 2 0 0 0 0 30 29 0 0 2
357 445
345 445
8 14 43 0 0 8320 0 30 35 0 0 4
363 427
285 427
285 529
266 529
6 13 44 0 0 8320 0 30 35 0 0 4
363 409
312 409
312 511
266 511
4 12 45 0 0 8320 0 30 35 0 0 4
363 391
303 391
303 493
266 493
2 11 46 0 0 8320 0 30 35 0 0 4
363 373
319 373
319 475
266 475
14 9 47 0 0 12416 0 34 30 0 0 4
265 376
291 376
291 436
363 436
7 13 48 0 0 4224 0 30 34 0 0 4
363 418
299 418
299 358
265 358
12 5 49 0 0 8320 0 34 30 0 0 4
265 340
308 340
308 400
363 400
3 11 50 0 0 8320 0 30 34 0 0 4
363 382
316 382
316 322
265 322
7 1 51 0 0 4224 0 40 32 0 0 4
150 157
47 157
47 153
48 153
6 0 2 0 0 0 0 40 0 0 112 4
150 148
145 148
145 188
137 188
0 0 2 0 0 0 0 0 0 115 113 2
137 179
137 206
8 0 2 0 0 0 0 40 0 0 114 5
150 166
137 166
137 206
136 206
136 223
1 0 2 0 0 0 0 33 0 0 0 4
137 241
137 223
136 223
136 219
2 5 2 0 0 0 0 40 40 0 0 6
150 112
137 112
137 179
137 179
137 139
150 139
2 1 2 0 0 0 0 40 40 0 0 4
150 112
150 147
150 147
150 103
8 4 52 0 0 12416 0 34 37 0 0 5
201 367
151 367
151 421
56 421
56 400
3 6 53 0 0 8320 0 37 34 0 0 5
62 400
62 413
158 413
158 349
201 349
2 4 54 0 0 8320 0 37 34 0 0 5
68 400
68 406
184 406
184 331
201 331
1 2 55 0 0 4224 0 37 34 0 0 4
74 400
168 400
168 313
201 313
9 4 56 0 0 12416 0 34 36 0 0 5
201 376
175 376
175 332
57 332
57 311
3 7 57 0 0 8320 0 36 34 0 0 5
63 311
63 328
180 328
180 358
201 358
5 2 58 0 0 4224 0 34 36 0 0 3
201 340
69 340
69 311
1 3 59 0 0 8320 0 36 34 0 0 3
75 311
75 322
201 322
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
