CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 270 30 130 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
110100498 256
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 389 515 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 Clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4460 0 0
2
42847.9 1
0
13 Logic Switch~
5 389 641 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 MODO
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3260 0 0
2
42847.9 0
0
9 Inverter~
13 657 522 0 2 22
0 19 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5156 0 0
2
42847.9 0
0
7 74LS190
134 711 549 0 14 29
0 21 20 17 18 12 11 10 9 35
36 23 24 25 26
0
0 0 4848 0
7 74LS190
-24 -51 25 -43
2 U1
-8 -52 6 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
3133 0 0
2
42847.9 0
0
12 Hex Display~
7 414 720 0 18 19
10 13 14 15 16 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5523 0 0
2
42847.9 1
0
12 Hex Display~
7 360 720 0 16 19
10 26 25 24 23 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3746 0 0
2
42847.9 0
0
7 74LS190
134 522 531 0 14 29
0 2 22 17 18 8 7 6 5 20
19 16 15 14 13
0
0 0 4848 0
7 74LS190
-24 -51 25 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 0 0 0 0 0
1 U
5668 0 0
2
42847.9 0
0
9 2-In AND~
219 1053 567 0 3 22
0 28 27 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5368 0 0
2
5.89797e-315 0
0
6 74LS85
106 922 362 0 14 29
0 23 24 25 26 2 2 3 2 32
33 34 28 37 38
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U2
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8293 0 0
2
5.89797e-315 5.36716e-315
0
6 74LS85
106 922 488 0 14 29
0 16 15 14 13 2 3 2 2 39
40 41 32 33 34
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3232 0 0
2
5.89797e-315 5.3568e-315
0
2 +V
167 823 299 0 1 3
0 3
0
0 0 53616 0
2 5V
-8 -22 6 -14
3 VCC
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6644 0 0
2
5.89797e-315 5.34643e-315
0
7 Ground~
168 859 839 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4978 0 0
2
5.89797e-315 5.32571e-315
0
6 74LS85
106 922 776 0 14 29
0 16 15 14 13 2 3 2 3 42
43 44 29 30 31
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9207 0 0
2
5.89797e-315 5.30499e-315
0
6 74LS85
106 922 650 0 14 29
0 23 24 25 26 2 2 2 2 29
30 31 45 46 27
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U6
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6998 0 0
2
5.89797e-315 5.26354e-315
0
7 74LS157
122 630 855 0 14 29
0 27 2 2 2 4 4 4 4 2
2 8 7 6 5
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3175 0 0
2
5.89797e-315 5.32571e-315
0
7 74LS157
122 630 738 0 14 29
0 27 2 2 2 2 4 2 2 2
2 12 11 10 9
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3378 0 0
2
5.89797e-315 5.30499e-315
0
2 +V
167 535 686 0 1 3
0 4
0
0 0 53616 0
2 5V
-8 -22 6 -14
4 VCC1
-13 -32 15 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
922 0 0
2
5.89797e-315 5.26354e-315
0
7 Ground~
168 562 920 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6891 0 0
2
5.89797e-315 0
0
7 Ground~
168 432 585 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5407 0 0
2
5.89797e-315 5.36716e-315
0
115
7 0 3 0 0 4096 0 9 0 0 100 2
890 389
823 389
8 0 2 0 0 4096 0 10 0 0 99 2
890 524
859 524
7 0 2 0 0 0 0 10 0 0 99 2
890 515
859 515
6 0 3 0 0 0 0 10 0 0 100 2
890 506
823 506
6 0 2 0 0 0 0 9 0 0 99 2
890 380
859 380
5 0 2 0 0 0 0 10 0 0 99 2
890 497
859 497
8 0 2 0 0 0 0 9 0 0 99 2
890 398
859 398
4 0 2 0 0 4096 0 15 0 0 110 2
598 846
562 846
8 0 2 0 0 0 0 16 0 0 110 2
598 765
562 765
6 0 4 0 0 4096 0 16 0 0 111 2
598 747
535 747
8 -143488 5 0 0 4096 0 7 0 0 113 2
490 567
451 567
7 -143487 6 0 0 4096 0 7 0 0 113 2
490 558
451 558
6 -143486 7 0 0 4096 0 7 0 0 113 2
490 549
451 549
5 -143485 8 0 0 4096 0 7 0 0 113 2
490 540
451 540
8 -143484 9 0 0 4096 0 4 0 0 112 2
679 585
649 585
7 -143483 10 0 0 4096 0 4 0 0 112 2
679 576
649 576
6 -143482 11 0 0 4096 0 4 0 0 112 2
679 567
649 567
5 -143481 12 0 0 4096 0 4 0 0 112 2
679 558
649 558
14 -656179328 13 0 0 4096 0 7 0 0 115 2
554 567
595 567
13 -656179327 14 0 0 4096 0 7 0 0 115 2
554 558
595 558
12 -656179326 15 0 0 4096 0 7 0 0 115 2
554 549
595 549
11 -656179325 16 0 0 4096 0 7 0 0 115 2
554 540
595 540
3 -13423565 17 0 0 4096 0 8 0 0 68 2
1074 567
1116 567
4 0 18 0 0 12416 0 4 0 0 25 4
679 549
620 549
620 641
414 641
4 1 18 0 0 0 0 7 2 0 0 4
490 531
414 531
414 641
401 641
10 1 19 0 0 4224 0 7 3 0 0 6
554 531
602 531
602 513
631 513
631 522
642 522
2 9 20 0 0 4224 0 4 7 0 0 4
679 531
612 531
612 522
560 522
2 1 21 0 0 4224 0 3 4 0 0 2
678 522
673 522
3 0 17 0 0 8192 0 7 0 0 62 3
484 522
465 522
465 469
2 1 22 0 0 4224 0 7 1 0 0 4
490 513
415 513
415 515
401 515
4 -656179321 23 0 0 4096 0 6 0 0 39 2
351 744
351 791
3 -656179322 24 0 0 4096 0 6 0 0 39 2
357 744
357 791
2 -656179323 25 0 0 4096 0 6 0 0 39 2
363 744
363 791
1 -656179324 26 0 0 4096 0 6 0 0 39 2
369 744
369 791
4 -656179325 16 0 0 4096 0 5 0 0 39 2
405 744
405 791
3 -656179326 15 0 0 4096 0 5 0 0 39 2
411 744
411 791
2 -656179327 14 0 0 4096 0 5 0 0 39 2
417 744
417 791
-656179328 1 13 0 0 4096 0 0 5 39 0 2
423 791
423 744
-160201 0 1 0 0 4128 0 0 0 0 0 2
450 791
324 791
1 0 2 0 0 0 0 7 0 0 114 2
484 504
475 504
-2475 0 1 0 0 32 0 0 0 0 0 2
432 436
432 488
1 0 27 0 0 4096 0 15 0 0 43 2
598 819
585 819
0 1 27 0 0 8320 0 0 16 63 0 5
1009 686
1009 919
585 919
585 702
598 702
8 0 4 0 0 0 0 15 0 0 111 2
598 882
535 882
6 0 4 0 0 0 0 15 0 0 111 2
598 864
535 864
2 0 2 0 0 0 0 15 0 0 110 2
598 828
562 828
4 0 2 0 0 0 0 16 0 0 110 2
598 729
562 729
2 0 2 0 0 0 0 16 0 0 110 2
598 711
562 711
10 0 2 0 0 0 0 16 0 0 110 2
592 783
562 783
10 0 2 0 0 0 0 15 0 0 110 2
592 900
562 900
9 0 2 0 0 0 0 15 0 0 110 2
598 891
562 891
7 0 4 0 0 0 0 15 0 0 111 2
598 873
535 873
5 0 4 0 0 0 0 15 0 0 111 2
598 855
535 855
3 0 2 0 0 0 0 15 0 0 110 2
598 837
562 837
9 0 2 0 0 0 0 16 0 0 110 2
598 774
562 774
7 0 2 0 0 0 0 16 0 0 110 2
598 756
562 756
5 0 2 0 0 0 0 16 0 0 110 2
598 738
562 738
3 0 2 0 0 0 0 16 0 0 110 2
598 720
562 720
8 0 3 0 0 0 0 13 0 0 100 2
890 812
823 812
7 0 2 0 0 0 0 13 0 0 99 2
890 803
859 803
6 0 3 0 0 0 0 13 0 0 100 2
890 794
823 794
-13423565 3 17 0 0 4224 0 0 4 41 0 4
432 469
621 469
621 540
673 540
14 2 27 0 0 0 0 14 8 0 0 4
954 686
1009 686
1009 576
1029 576
14 -656179324 26 0 0 0 0 4 0 0 98 2
743 585
783 585
13 -656179323 25 0 0 0 0 4 0 0 98 2
743 576
783 576
12 -656179322 24 0 0 0 0 4 0 0 98 2
743 567
783 567
11 -656179321 23 0 0 0 0 4 0 0 98 2
743 558
783 558
-2475 0 1 0 0 48 0 0 0 0 0 2
1116 535
1116 587
12 1 28 0 0 8320 0 9 8 0 0 4
954 380
1009 380
1009 558
1029 558
5 0 2 0 0 0 0 13 0 0 99 2
890 785
859 785
8 0 2 0 0 0 0 14 0 0 99 2
890 686
859 686
5 0 2 0 0 0 0 14 0 0 99 2
890 659
859 659
6 0 2 0 0 0 0 14 0 0 99 2
890 668
859 668
7 0 2 0 0 0 0 14 0 0 99 2
890 677
859 677
4 -656179328 13 0 0 4224 0 13 0 0 98 2
890 776
783 776
3 -656179327 14 0 0 4224 0 13 0 0 98 2
890 767
783 767
2 -656179326 15 0 0 4224 0 13 0 0 98 2
890 758
783 758
1 -656179325 16 0 0 4224 0 13 0 0 98 2
890 749
783 749
4 -656179324 26 0 0 4224 0 14 0 0 98 2
890 650
783 650
3 -656179323 25 0 0 4224 0 14 0 0 98 2
890 641
783 641
2 -656179322 24 0 0 4224 0 14 0 0 98 2
890 632
783 632
1 -656179321 23 0 0 4224 0 14 0 0 98 2
890 623
783 623
9 12 29 0 0 8320 0 14 13 0 0 4
954 623
985 623
985 794
954 794
13 10 30 0 0 8320 0 13 14 0 0 4
954 803
976 803
976 632
954 632
14 11 31 0 0 8320 0 13 14 0 0 4
954 812
968 812
968 641
954 641
3 -656179327 14 0 0 0 0 10 0 0 98 2
890 479
783 479
2 -656179326 15 0 0 0 0 10 0 0 98 2
890 470
783 470
1 -656179325 16 0 0 0 0 10 0 0 98 2
890 461
783 461
3 -656179323 25 0 0 0 0 9 0 0 98 2
890 353
783 353
2 -656179322 24 0 0 0 0 9 0 0 98 2
890 344
783 344
1 -656179321 23 0 0 0 0 9 0 0 98 2
890 335
783 335
5 0 2 0 0 0 0 9 0 0 99 2
890 371
859 371
4 -656179328 13 0 0 0 0 10 0 0 98 2
890 488
783 488
4 -656179324 26 0 0 0 0 9 0 0 98 2
890 362
783 362
9 12 32 0 0 8320 0 9 10 0 0 4
954 335
985 335
985 506
954 506
13 10 33 0 0 8320 0 10 9 0 0 4
954 515
976 515
976 344
954 344
14 11 34 0 0 8320 0 10 9 0 0 4
954 524
968 524
968 353
954 353
-160201 0 1 0 0 4256 0 0 0 0 0 2
783 290
783 851
1 0 2 0 0 4224 0 12 0 0 0 2
859 833
859 298
1 0 3 0 0 4224 0 11 0 0 0 2
823 308
823 848
14 -143488 5 0 0 4224 0 15 0 0 109 2
662 891
721 891
13 -143487 6 0 0 4224 0 15 0 0 109 2
662 873
721 873
12 -143486 7 0 0 4224 0 15 0 0 109 2
662 855
721 855
11 -143485 8 0 0 4224 0 15 0 0 109 2
662 837
721 837
14 -143484 9 0 0 4224 0 16 0 0 109 2
662 774
721 774
13 -143483 10 0 0 4224 0 16 0 0 109 2
662 756
721 756
12 -143482 11 0 0 4224 0 16 0 0 109 2
662 738
721 738
11 -143481 12 0 0 4224 0 16 0 0 109 2
662 720
721 720
-144841 0 1 0 0 32 0 0 0 0 0 2
721 683
721 911
1 0 2 0 0 0 0 18 0 0 0 2
562 914
562 684
1 0 4 0 0 4224 0 17 0 0 0 2
535 695
535 919
-144841 0 1 0 0 32 0 0 0 0 0 2
649 627
649 553
-144841 0 1 0 0 32 0 0 0 0 0 2
451 611
451 536
0 1 2 0 0 0 0 0 19 0 0 3
485 504
432 504
432 579
-160201 0 1 0 0 32 0 0 0 0 0 2
595 631
595 535
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
