CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 920 30 80 10
176 80 1278 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
57
13 Logic Switch~
5 124 1502 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 A14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8132 0 0
2
42814.5 4
0
13 Logic Switch~
5 122 1420 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 A13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
65 0 0
2
42814.5 3
0
13 Logic Switch~
5 124 1339 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 A12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6609 0 0
2
42814.5 2
0
13 Logic Switch~
5 126 1259 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 A11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8995 0 0
2
42814.5 1
0
13 Logic Switch~
5 125 1172 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 A10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3918 0 0
2
42814.5 0
0
13 Logic Switch~
5 139 678 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7519 0 0
2
42814.5 4
0
13 Logic Switch~
5 140 765 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
377 0 0
2
42814.5 3
0
13 Logic Switch~
5 138 845 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8816 0 0
2
42814.5 2
0
13 Logic Switch~
5 136 926 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3877 0 0
2
42814.5 1
0
13 Logic Switch~
5 138 1008 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
926 0 0
2
42814.5 0
0
13 Logic Switch~
5 135 524 0 1 11
0 47
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7262 0 0
2
5.89793e-315 5.26354e-315
0
13 Logic Switch~
5 133 442 0 1 11
0 49
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5267 0 0
2
5.89793e-315 5.26354e-315
0
13 Logic Switch~
5 135 361 0 1 11
0 52
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8838 0 0
2
5.89793e-315 5.26354e-315
0
13 Logic Switch~
5 137 281 0 1 11
0 50
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7159 0 0
2
5.89793e-315 5.26354e-315
0
13 Logic Switch~
5 136 194 0 1 11
0 55
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5812 0 0
2
5.89793e-315 0
0
10 8-In NAND~
219 1170 1365 0 9 19
0 6 5 4 3 2 2 2 2 7
0
0 0 624 0
6 74LS30
-21 -24 21 -16
2 U3
-8 -44 6 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 0 0 0 0
1 U
331 0 0
2
42814.6 0
0
9 Inverter~
13 205 1500 0 2 22
0 10 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not2C
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 15 0
1 U
9604 0 0
2
42814.5 19
0
9 Inverter~
13 203 1418 0 2 22
0 11 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not2B
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 15 0
1 U
7518 0 0
2
42814.5 18
0
9 Inverter~
13 205 1337 0 2 22
0 14 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not2A
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 15 0
1 U
4832 0 0
2
42814.5 17
0
9 Inverter~
13 207 1257 0 2 22
0 12 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not1F
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
6798 0 0
2
42814.5 16
0
9 Inverter~
13 206 1170 0 2 22
0 17 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not1E
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
3336 0 0
2
42814.5 15
0
14 Logic Display~
6 1270 1222 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8370 0 0
2
42814.5 14
0
5 7422~
219 872 1478 0 5 22
0 15 8 14 10 2
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U8B
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 13 0
1 U
3910 0 0
2
42814.5 13
0
5 7412~
219 768 1400 0 4 22
0 17 13 9 3
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 14 0
1 U
316 0 0
2
42814.5 12
0
5 7412~
219 779 1328 0 4 22
0 17 12 11 4
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 14 0
1 U
536 0 0
2
42814.5 11
0
5 7412~
219 787 1237 0 4 22
0 12 13 9 5
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 14 0
1 U
4460 0 0
2
42814.5 10
0
5 7422~
219 788 1100 0 5 22
0 16 14 15 8 6
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U8A
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 13 0
1 U
3260 0 0
2
42814.5 9
0
10 2-In NAND~
219 1195 984 0 3 22
0 19 18 27
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
5156 0 0
2
42814.5 0
0
10 2-In NAND~
219 1073 755 0 3 22
0 21 20 19
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3133 0 0
2
42814.5 0
0
10 2-In NAND~
219 934 865 0 3 22
0 25 26 20
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5523 0 0
2
42814.5 0
0
10 2-In NAND~
219 939 675 0 3 22
0 23 24 21
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3746 0 0
2
42814.5 0
0
5 7422~
219 804 641 0 5 22
0 35 33 34 22 23
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U4B
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 11 0
1 U
5668 0 0
2
42814.5 0
0
5 7412~
219 804 734 0 4 22
0 31 32 28 24
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 12 0
1 U
5368 0 0
2
42814.5 0
0
5 7412~
219 800 827 0 4 22
0 36 31 30 25
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 12 0
1 U
8293 0 0
2
42814.5 0
0
5 7412~
219 800 930 0 4 22
0 36 32 28 26
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 12 0
1 U
3232 0 0
2
42814.5 0
0
5 7422~
219 791 1025 0 5 22
0 34 22 33 29 18
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U4A
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 11 0
1 U
6644 0 0
2
42814.5 0
0
14 Logic Display~
6 1284 728 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4978 0 0
2
42814.5 19
0
9 Inverter~
13 220 676 0 2 22
0 36 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not1D
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
9207 0 0
2
42814.5 18
0
9 Inverter~
13 221 763 0 2 22
0 31 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not1C
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
6998 0 0
2
42814.5 17
0
9 Inverter~
13 219 843 0 2 22
0 33 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not1B
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
3175 0 0
2
42814.5 16
0
9 Inverter~
13 217 924 0 2 22
0 30 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
5 Not1A
-17 -29 18 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
3378 0 0
2
42814.5 15
0
9 Inverter~
13 219 1006 0 2 22
0 29 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotF
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
922 0 0
2
42814.5 14
0
8 2-In OR~
219 1189 500 0 3 22
0 42 37 41
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
6891 0 0
2
5.89793e-315 0
0
8 2-In OR~
219 1051 271 0 3 22
0 43 38 42
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
5407 0 0
2
5.89793e-315 0
0
8 2-In OR~
219 934 382 0 3 22
0 40 39 38
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
7349 0 0
2
5.89793e-315 0
0
8 2-In OR~
219 925 191 0 3 22
0 45 44 43
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3919 0 0
2
5.89793e-315 0
0
9 3-In AND~
219 799 445 0 4 22
0 55 51 46 39
0
0 0 624 0
5 74F11
-18 -28 17 -20
5 Caso4
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 4 0
1 U
9747 0 0
2
5.89793e-315 5.34643e-315
0
9 3-In AND~
219 798 343 0 4 22
0 55 50 49 40
0
0 0 624 0
5 74F11
-18 -28 17 -20
5 Caso3
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 4 0
1 U
5310 0 0
2
5.89793e-315 5.32571e-315
0
9 3-In AND~
219 798 250 0 4 22
0 50 51 46 44
0
0 0 624 0
5 74F11
-18 -28 17 -20
5 Caso2
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
4318 0 0
2
5.89793e-315 5.30499e-315
0
9 4-In AND~
219 798 156 0 5 22
0 54 53 52 48 45
0
0 0 624 0
6 74LS21
-21 -28 21 -20
5 Caso1
-19 -28 16 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
3917 0 0
2
5.89793e-315 5.26354e-315
0
9 4-In AND~
219 801 544 0 5 22
0 53 52 48 47 37
0
0 0 624 0
6 74LS21
-21 -28 21 -20
5 Caso5
-19 -28 16 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
7930 0 0
2
5.89793e-315 0
0
9 Inverter~
13 216 522 0 2 22
0 47 46
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotE
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
6128 0 0
2
5.89793e-315 0
0
9 Inverter~
13 214 440 0 2 22
0 49 48
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotD
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
7346 0 0
2
5.89793e-315 0
0
9 Inverter~
13 216 359 0 2 22
0 52 51
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotC
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8577 0 0
2
5.89793e-315 0
0
9 Inverter~
13 218 279 0 2 22
0 50 53
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotB
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3372 0 0
2
5.89793e-315 0
0
9 Inverter~
13 217 192 0 2 22
0 55 54
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotA
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3741 0 0
2
5.89793e-315 5.26354e-315
0
14 Logic Display~
6 1281 244 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5813 0 0
2
5.89793e-315 0
0
107
8 0 2 0 0 8192 0 16 0 0 4 3
1146 1397
1146 1398
1115 1398
7 0 2 0 0 0 0 16 0 0 4 3
1146 1388
1146 1389
1115 1389
6 0 2 0 0 0 0 16 0 0 4 3
1146 1379
1146 1380
1115 1380
5 5 2 0 0 4224 0 23 16 0 0 5
899 1478
1115 1478
1115 1371
1146 1371
1146 1370
4 4 3 0 0 8320 0 16 24 0 0 5
1146 1361
1146 1362
854 1362
854 1400
795 1400
4 3 4 0 0 4224 0 25 16 0 0 5
806 1328
1079 1328
1079 1353
1146 1353
1146 1352
4 2 5 0 0 4224 0 26 16 0 0 5
814 1237
1090 1237
1090 1344
1146 1344
1146 1343
5 1 6 0 0 4224 0 27 16 0 0 5
815 1100
1102 1100
1102 1335
1146 1335
1146 1334
9 1 7 0 0 12416 0 16 22 0 0 4
1197 1365
1197 1366
1270 1366
1270 1240
2 0 8 0 0 8192 0 23 0 0 14 5
848 1484
802 1484
802 1583
761 1583
761 1610
0 3 9 0 0 4096 0 0 26 12 0 4
635 1433
620 1433
620 1246
763 1246
2 3 9 0 0 4224 0 17 24 0 0 4
226 1500
635 1500
635 1409
744 1409
4 0 10 0 0 20608 0 23 0 0 28 7
848 1496
821 1496
821 1536
591 1536
591 1458
143 1458
143 1500
0 0 8 0 0 8208 0 0 0 15 0 3
549 1418
549 1610
766 1610
2 4 8 0 0 4224 0 18 27 0 0 7
224 1418
549 1418
549 1181
762 1181
762 1145
764 1145
764 1118
3 0 11 0 0 12416 0 25 0 0 29 5
755 1337
508 1337
508 1374
143 1374
143 1418
0 0 12 0 0 4096 0 0 0 24 31 3
371 1219
138 1219
138 1257
0 2 13 0 0 8192 0 0 24 19 0 3
472 1337
472 1400
744 1400
2 2 13 0 0 12416 0 19 26 0 0 4
226 1337
472 1337
472 1237
763 1237
0 3 14 0 0 8192 0 0 23 21 0 3
437 1288
437 1472
848 1472
0 2 14 0 0 8320 0 0 27 30 0 7
143 1337
143 1288
437 1288
437 1139
715 1139
715 1106
764 1106
0 1 15 0 0 8192 0 0 23 23 0 4
403 1257
403 1452
848 1452
848 1460
2 3 15 0 0 12416 0 20 27 0 0 4
228 1257
403 1257
403 1094
764 1094
1 2 12 0 0 4224 0 26 25 0 0 6
763 1228
371 1228
371 1219
371 1219
371 1328
755 1328
2 1 16 0 0 12416 0 21 27 0 0 5
227 1170
341 1170
341 1077
764 1077
764 1082
0 1 17 0 0 8320 0 0 24 27 0 3
287 1312
287 1391
744 1391
0 1 17 0 0 0 0 0 25 32 0 5
139 1172
139 1126
287 1126
287 1319
755 1319
1 1 10 0 0 0 0 1 17 0 0 3
136 1502
136 1500
190 1500
1 1 11 0 0 0 0 2 18 0 0 3
134 1420
134 1418
188 1418
1 1 14 0 0 0 0 3 19 0 0 3
136 1339
136 1337
190 1337
1 1 12 0 0 0 0 4 20 0 0 3
138 1259
138 1257
192 1257
1 1 17 0 0 0 0 5 21 0 0 4
137 1172
139 1172
139 1170
191 1170
2 0 18 0 0 4096 0 28 0 0 46 2
1171 993
1174 993
1 0 19 0 0 4096 0 28 0 0 51 2
1171 975
1174 975
2 0 20 0 0 4096 0 29 0 0 47 2
1049 764
1037 764
1 0 21 0 0 4096 0 29 0 0 52 2
1049 746
1037 746
3 0 20 0 0 0 0 30 0 0 47 3
961 865
961 866
973 866
3 0 21 0 0 0 0 31 0 0 52 2
966 675
966 675
4 0 22 0 0 4096 0 32 0 0 59 3
780 659
780 654
775 654
5 0 23 0 0 8192 0 32 0 0 54 4
831 641
831 639
826 639
826 640
4 0 24 0 0 4096 0 33 0 0 53 2
831 734
828 734
4 0 25 0 0 0 0 34 0 0 49 2
827 827
827 827
4 0 26 0 0 4096 0 35 0 0 48 2
827 930
827 929
2 0 22 0 0 8192 0 36 0 0 58 3
767 1031
767 1033
775 1033
5 0 18 0 0 8192 0 36 0 0 46 4
818 1025
818 1029
830 1029
830 1028
0 0 18 0 0 4224 0 0 0 0 0 4
825 1028
1125 1028
1125 993
1179 993
0 0 20 0 0 8320 0 0 0 0 0 4
970 866
1009 866
1009 764
1041 764
2 0 26 0 0 12416 0 30 0 0 0 5
910 874
910 875
869 875
869 929
823 929
0 1 25 0 0 4224 0 0 30 0 0 5
822 827
869 827
869 857
910 857
910 856
3 1 27 0 0 8320 0 28 37 0 0 3
1222 984
1284 984
1284 746
3 0 19 0 0 8320 0 29 0 0 0 4
1100 755
1125 755
1125 975
1179 975
0 0 21 0 0 8320 0 0 0 0 0 4
961 675
1009 675
1009 746
1041 746
2 0 24 0 0 8320 0 31 0 0 0 4
915 684
869 684
869 734
822 734
0 1 23 0 0 4224 0 0 31 0 0 4
822 640
869 640
869 666
915 666
0 3 28 0 0 4096 0 0 33 56 0 3
634 939
634 743
780 743
2 3 28 0 0 4224 0 42 35 0 0 4
240 1006
634 1006
634 939
776 939
4 0 29 0 0 16512 0 36 0 0 72 6
767 1043
767 1042
605 1042
605 964
157 964
157 1006
0 0 22 0 0 8192 0 0 0 59 0 3
563 924
563 1033
780 1033
2 0 22 0 0 4224 0 41 0 0 0 5
238 924
563 924
563 654
776 654
776 651
3 0 30 0 0 12416 0 34 0 0 73 5
776 836
522 836
522 880
157 880
157 924
0 0 31 0 0 4096 0 0 0 68 75 3
385 725
152 725
152 763
0 2 32 0 0 8192 0 0 35 63 0 3
486 843
486 930
776 930
2 2 32 0 0 12416 0 40 33 0 0 4
240 843
486 843
486 734
780 734
0 3 33 0 0 8192 0 0 36 65 0 3
451 794
451 1019
767 1019
0 2 33 0 0 16512 0 0 32 74 0 6
157 843
157 794
451 794
451 645
780 645
780 647
0 1 34 0 0 8192 0 0 36 67 0 4
417 763
417 1015
767 1015
767 1007
2 3 34 0 0 12416 0 39 32 0 0 4
242 763
417 763
417 635
780 635
1 2 31 0 0 4224 0 33 34 0 0 4
780 725
385 725
385 827
776 827
2 1 35 0 0 12416 0 38 32 0 0 5
241 676
355 676
355 627
780 627
780 623
0 1 36 0 0 8320 0 0 35 71 0 3
301 818
301 921
776 921
0 1 36 0 0 0 0 0 34 76 0 5
153 678
153 632
301 632
301 818
776 818
1 1 29 0 0 0 0 10 42 0 0 3
150 1008
150 1006
204 1006
1 1 30 0 0 0 0 9 41 0 0 3
148 926
148 924
202 924
1 1 33 0 0 0 0 8 40 0 0 3
150 845
150 843
204 843
1 1 31 0 0 0 0 7 39 0 0 3
152 765
152 763
206 763
1 1 36 0 0 0 0 6 38 0 0 4
151 678
153 678
153 676
205 676
5 2 37 0 0 4224 0 51 43 0 0 4
822 544
1122 544
1122 509
1176 509
3 2 38 0 0 8320 0 45 44 0 0 4
967 382
1006 382
1006 280
1038 280
2 4 39 0 0 4224 0 45 47 0 0 4
921 391
866 391
866 445
820 445
4 1 40 0 0 12416 0 48 45 0 0 4
819 343
866 343
866 373
921 373
3 1 41 0 0 8320 0 43 57 0 0 3
1222 500
1281 500
1281 262
3 1 42 0 0 8320 0 44 43 0 0 4
1084 271
1122 271
1122 491
1176 491
3 1 43 0 0 8320 0 46 44 0 0 4
958 191
1006 191
1006 262
1038 262
2 4 44 0 0 8320 0 46 49 0 0 4
912 200
866 200
866 250
819 250
5 1 45 0 0 4224 0 50 46 0 0 4
819 156
866 156
866 182
912 182
0 3 46 0 0 4096 0 0 49 87 0 3
631 455
631 259
774 259
2 3 46 0 0 4224 0 52 47 0 0 4
237 522
631 522
631 454
775 454
4 0 47 0 0 12416 0 51 0 0 103 5
777 558
602 558
602 480
154 480
154 522
0 3 48 0 0 8192 0 0 51 90 0 3
560 440
560 549
777 549
2 4 48 0 0 4224 0 53 50 0 0 4
235 440
560 440
560 170
774 170
3 0 49 0 0 12416 0 48 0 0 104 5
774 352
519 352
519 396
154 396
154 440
0 0 50 0 0 4096 0 0 0 99 106 3
382 241
149 241
149 279
0 2 51 0 0 8320 0 0 47 94 0 3
483 359
483 445
775 445
2 2 51 0 0 0 0 54 49 0 0 4
237 359
483 359
483 250
774 250
0 2 52 0 0 8320 0 0 51 96 0 3
448 310
448 540
777 540
0 3 52 0 0 0 0 0 50 105 0 5
154 359
154 310
448 310
448 161
774 161
0 1 53 0 0 8320 0 0 51 98 0 3
414 279
414 531
777 531
2 2 53 0 0 0 0 55 50 0 0 4
239 279
414 279
414 152
774 152
1 2 50 0 0 4224 0 49 48 0 0 4
774 241
382 241
382 343
774 343
2 1 54 0 0 12416 0 56 50 0 0 4
238 192
352 192
352 143
774 143
0 1 55 0 0 8320 0 0 47 102 0 3
298 334
298 436
775 436
0 1 55 0 0 0 0 0 48 107 0 5
150 194
150 148
298 148
298 334
774 334
1 1 47 0 0 0 0 11 52 0 0 3
147 524
147 522
201 522
1 1 49 0 0 0 0 12 53 0 0 3
145 442
145 440
199 440
1 1 52 0 0 0 0 13 54 0 0 3
147 361
147 359
201 359
1 1 50 0 0 0 0 14 55 0 0 3
149 281
149 279
203 279
1 1 55 0 0 0 0 15 56 0 0 4
148 194
150 194
150 192
202 192
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
